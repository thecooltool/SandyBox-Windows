MZP      ��  �       @    �!jr                             � �	�!�L�!��This program must be run under Win32
$7                                                                                                                                                                                                                                                                                                                                                                                                        PE  L %ӖS        � #                         @                      �                                                    �                                                                                                         .text                                `.data                             @  �.rsrc    �     �                @  @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    a]�D          @  �   `  �   �  �
   X �   � �   � �    a]�D          � �   � �    a]�D       y   �y    �y  8 �    a]�D      x    P �   h �   � �   � �	   � �
   � �   � �   � �    �   ( �   @ �   X �   p �   � �   � �   � �   � �   � �     �    �   0 �   H �   ` �   x �   � �    � �!   � �"   � �&   � �'   	 �(    	 �,   8	 �B   P	 �E   h	 �F   �	 �G   �	 �H   �	 �I   �	 �J   �	 �R   �	 �S   
 �T   (
 �U   @
 �V   X
 �X   p
 �Y   �
 �\   �
 �]   �
 �^   �
 �_   �
 �`     �e    �f   0 �g   H �h   ` �i   x �j   � �k   � �l   � �m   � �n   � �o    �p     �q   8 �r   P �s   h �t   � �u   � �w   � �x   � �~   � �   � ��    ��   ( ��   @ ��   X ��   p ��   � ��   � �  � �  � �  � �    �   �  0 �  H �  ` ��  x ��  � ��  � ��  � ��  � ��  � ��   ��    ��  8 ��  P ��  h ��  � ��  � ��  � ��  � ��  � ��  � ��   ��  ( ��  @ ��  X ��  p ��  � ��  � ��  � ��  � ��  � ��    ��   ��  0 ��  H ��  ` �   x �    a]�D    (   � �� �� �� �  �� �<  �� �Z  �� �x  � ��  �  ��  �8 ��  �P �! �h �<! �� �f! �� ��! �� ��! �� ��! �� ��! �� �" � �:" �( �f" �@ ��" �X ��" �p ��" �� �# �� � # �� �:# �� �d# �� ��# �  ��# � ��# �0 ��# �H � $ �` �@$ �x �Z$ �� �~$ �� ��$ �� ��$ �� ��$ �� �
% � �B% �  �h% �8 �    a]�D       y  P �    a]�D          h �    a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D                a]�D               a]�D                a]�D         0      a]�D         @      a]�D         P      a]�D         `      a]�D         p      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D                a]�D               a]�D                a]�D         0      a]�D         @      a]�D         P      a]�D         `      a]�D         p      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D                a]�D               a]�D                a]�D         0      a]�D         @      a]�D         P      a]�D         `      a]�D         p      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D                a]�D               a]�D                a]�D         0      a]�D         @      a]�D         P      a]�D         `      a]�D         p      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D                a]�D               a]�D                a]�D         0      a]�D         @      a]�D         P      a]�D         `      a]�D         p      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D                a]�D               a]�D                a]�D         0      a]�D         @      a]�D         P      a]�D         `      a]�D         p      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D                a]�D               a]�D                a]�D         0      a]�D         @      a]�D         P      a]�D         `      a]�D         p      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D         �      a]�D                a]�D               a]�D                a]�D         0      a]�D         @      a]�D           P      a]�D           `      a]�D           p      a]�D           �      a]�D           �      a]�D           �      a]�D           �      a]�D           �      a]�D           �      a]�D           �      a]�D           �      a]�D                  a]�D                 a]�D                  a]�D           0      a]�D           @      a]�D           P      a]�D           `      a]�D           p      a]�D           �      a]�D           �      a]�D           �      a]�D           �      a]�D           �      a]�D           �      a]�D           �      a]�D           �      a]�D                  a]�D                 a]�D                  a]�D           0      a]�D           @      a]�D           P      a]�D           `      a]�D           p      a]�D           �      a]�D           �      a]�D           �      a]�D           �      a]�D           �      a]�D         �      a]�D         �  �5  4          �6  �           �7  �           <8  l          �9  D          �:  �!          |\  �D          L�  J          ��  l          �            $�  v          ��  �          ��  ^          ��  �          ��  �          h�            p�  :          ��  �          |�  &          ��  T          ��  p          h�  �          �  �          �  �           ��  J          �  �          � P          � &           �            �          � r          \           t �            �          � �          x �             D          \! �          L7 �            8 d          �; 2          �C           �Q �          PY *          |\           �c h          �g V          L} �          � �          Ԏ �          p� �          � .          4�           H� 8          �� �          H� �          @� z          �� F          � n          t� v           � *          � �          Ժ �          �� �          P� �          � �          �� �          �� �          \�           t� �          $� "          H� N          �� X          �� F          8�           H�           `�            `� Z          �� p          ,� (          T� l           �� �           �� �           �           0� >           p� J          �� �          H� �          �� �          �� �           t� �          8 d          �           � \           �          � �          T �          � 4          " �          % t          �& �           L' �          ) 
           - �          �0 �          �3 D          $8 �          �: z          p> �          pE `          �I h          8M           XP j          �T R          Y            8] �          �` v          hc �          dg $          �h �           |i �          @l            `n v          �q            �u �          �y            �y ο         �9 [          �F �          �M P6          � Ph          h� �          �� �
          �� O          0 �          � l
          D �          �  R          P9 ^          �D U�           �
          �' �          �;           �K �          $c �          �i ]          Pl �B          � �          �� ~�           I Y�          |7 ^          �L &�           	 -          4.	 �          �B	 �          `N	 `          �R	 o[          0�	 �          42
 T          P�
           `�
 ͗          0$ �           * �z          � P          0� �          �� "           �� D           D V C L A L  T A B O U T D I A L O G  T A U T H E N T I C A T E F O R M  T C L E A N U P D I A L O G  T C O N S O L E D I A L O G  T C O P Y D I A L O G  T C O P Y P A R A M C U S T O M D I A L O G  T C O P Y P A R A M P R E S E T D I A L O G  T C O P Y P A R A M S F R A M E  T C R E A T E D I R E C T O R Y D I A L O G  T C U S T O M C O M M A N D D I A L O G  T C U S T O M D I A L O G  T C U S T O M S C P E X P L O R E R F O R M  T E D I T M A S K D I A L O G  T E D I T O R F O R M  T E D I T O R P R E F E R E N C E S D I A L O G  T F I L E F I N D D I A L O G  T F I L E S Y S T E M I N F O D I A L O G  T F U L L S Y N C H R O N I Z E D I A L O G  T I M P O R T S E S S I O N S D I A L O G  T L I C E N S E D I A L O G  T L O C A T I O N P R O F I L E S D I A L O G  T L O G F O R M  T L O G I N D I A L O G  T N O N V I S U A L D A T A M O D U L E  T O P E N D I R E C T O R Y D I A L O G  T P R E F E R E N C E S D I A L O G  T P R O G R E S S F O R M  T P R O P E R T I E S D I A L O G  T R E M O T E T R A N S F E R D I A L O G  T R I G H T S E X T F R A M E  T R I G H T S F R A M E  T S C P C O M M A N D E R F O R M  T S C P E X P L O R E R F O R M  T S E L E C T M A S K D I A L O G  T S I T E A D V A N C E D D I A L O G  T S Y M L I N K D I A L O G  T S Y N C H R O N I Z E C H E C K L I S T D I A L O G  T S Y N C H R O N I Z E D I A L O G  T S Y N C H R O N I Z E P R O G R E S S F O R M     (       @                                ���                                  8   0   p   `   �   �  �  �  �  �  �  �  �  �  �                                 ����������������������������������������������������?��?��?� �?�  ?�  �p ���������������������������  (                �                       ��� �  �  ��  �H  �x  �H  ��  �d  ��  �)  �9  �  ��  �|  �   �   �  �  x  0�  �  �         !              �  �  ?�  (      
         P                         �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ��� �����  �����  �www�  �  �  ����  �  �  �����  �����  �����          (   '                                    �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                     ����� ����  ����� ����� ������ ����� ���� ����� ����� ������ ����� ���� ����� ����� ������ ����� ���� ����� ����� ������ ����� ���� ����� ����� ������ ����� ����  �����                     (   !            �                         �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ��� �����������������   ������������wwww�   ������������w�ww�   ������� ���x�ww�   �������  ������w�   ������� ���x�w�   ��������� ���w���   ��������� ��wwx��   ������������www��   ������������wwww�   �����������������     �* * F o r t s � t t   a n s l u t a   t i l l   e n   o k � n d   s e r v e r   o c h   l � g g a   t i l l   d e s s   v � r d n y c k e l   t i l l   c a c h e n ? * * 
 
 S e r v e r n s   v � r d n y c k e l   h i t t a d e s   i n t e   i   c a c h e n .   D u   h a r   i n g e n   g a r a n t i   a t t   s e r v e r n   � r   d e n   d a t o r   s o m   d u   t r o r   a t t   d e t   � r . 
 
 S e r v e r n s   % s   f i n g e r a v t r y c k s n y c k e l   � r : 
 % s 
 O m   d u   l i t a r   p �   d e n n a   v � r d ,   t r y c k   p �   J a .   F � r   a t t   a n s l u t a   u t a n   a t t   v � r d n y c k e l n   l � g g s   t i l l   c a c h e n ,   t r y c k   p �   N e j .   F � r   a t t   a v b r y t a   a n s l u t n i n g e n   t r y c k   p �   A v b r y t .  * * V A R N I N G   -   S � K E R H E T S R I S K ! * * 
 
 S e r v e r n s   v � r d n y c k e l   m a t c h a r   i n t e   d e n   s o m   W i n S C P   h a r   i   c a c h e n .   D e t   i n n e b � r   a t t   a n t i n g e n   s e r v e r a d m i n i s t r a t � r e n   h a r   � n d r a t   v � r d n y c k e l n   ( s e r v e r n   p r e s e n t e r a r   o l i k a   n y c k l a r   u n d e r   v i s s a   o m s t � n d i g h e t e r )   e l l e r   a t t   d u   h a r   a n s l u t i t   t i l l   e n   a n n a n   d a t o r   s o m   l � t s a s   v a r a   s e r v e r n . 
 
 D e n   n y a   % s   f i n g e r a v t r y c k s n y c k e l n   � r : 
 % s 
 
 O m   d u   v � n t a d e   d e n n a   f � r � n d r i n g ,   l i t a r   p �   d e n   n y a   n y c k e l n   o c h   v i l l   f o r t s � t t a   a t t   a n s l u t a   t i l l   s e r v e r n ,   a n t i n g e n   t r y c k   p �   ' U p p d a t e r a '   f � r   a t t   u p p d a t e r a   c a c h e n   e l l e r   t r y c k   p �   ' L � g g   t i l l '   f � r   a t t   l � g g a   t i l l   d e n   n y a   n y c k e l n   i   c a c h e n   s a m t i d i g t   s o m   d e n   g a m l a   b e h � l l s .   O m   d u   v i l l   f o r t s � t t a   a n s l u t a ,   m e n   u t a n   a t t   u p p d a t e r a   c a c h e n ,   t r y c k   p �   ' H o p p a   � v e r ' .   O m   d u   v i l l   a v b r y t a   a n s l u t n i n g e n   h e l t   t r y c k e r   d u   p �   ' A v b r y t ' .   A t t   t r y c k a   p �   A v b r y t   � r   d e t   E N D A   g a r a n t e r a t   s � k r a   v a l e t . 0D u   l a d d a r   e n   S S H - 2   p r i v a t   n y c k e l   s o m   h a r   e t t   g a m m a l t   f i l f o r m a t .   D e t   i n n e b � r   a t t   d i n   n y c k e l f i l   i n t e   � r   h e l t   s � k e r   f � r   m a n i p u l e r i n g s f � r s � k .   V i   r e k o m m e n d e r a r   d i g   a t t   k o n v e r t e r a   d i n   n y c k e l   t i l l   d e t   n y a   f o r m a t e t . 
 
 D u   k a n   u t f � r a   d e n   h � r   k o n v e r t e r i n g e n   g e n o m   a t t   l a d d a   f i l e n   i   P u T T Y g e n   o c h   s e d a n   s p a r a   d e n   i g e n . � H e l p   [   < k o m m a n d o >   [   < k o m m a n d o 2 >   . . .   ] 
     V i s a r   l i s t a   p �   k o m m a n d o n   o m   i n g a   p a r a m e t e r a r   a n g e s . 
     V i s a r   h j � l p   o m   e t t   k o m m a n d o   o m   d e t   a n g e s . 
 a l i a s : 
     m a n 
 e x e m p e l : 
     h e l p 
     h e l p   l s 
 D e x i t 
     S t � n g e r   a l l a   s e s s i o n e r   o c h   a v s l u t a r   p r o g r a m m e t . 
 a l i a s : 
     b y e 
 �o p e n   < w e b b p l a t s > 
 o p e n   [   s f t p | s c p | f t p : / /   ] [ < a n v � n d a r e >   [   : l � s e n o r d   ]   @   ]   < v � r d >   [   : < p o r t > 
   U p p r � t t a r   a n s l u t n i n g   t i l l   g i v e n   v � r d .   A n v � n d   a n t i n g e n   n a m n e t   p �   w e b b p l a t s e n   e l l e r 
   n a m n g e   v � r d ,   a n v � n d a r n a m n ,   p o r t ,   o c h   p r o t o k o l l   d i r e k t . 
 v � x l a r : 
   - p r i v a t e k e y = < n y c k e l >     P r i v a t   n y c k e l f i l 
     - t i m e o u t = < s e k >           T i m e o u t   f � r   s e r v e r s v a r 
     - h o s t k e y = < f i n g e r a v t r y c k >   F i n g e r a v t r y c k   f � r   s e r v e r n   v � r d n y c k e l   ( e n d a s t   S F T P   o c h   S C P ) . 
     - c e r t i f i c a t e = < f i n g e r a v t r y c k >   F i n g e r a v t r y c k   f � r   S S L / T L S   c e r t i f i k a t   ( e n d a s t   F T P S ) 
     - p a s s i v e = o n | o f f         P a s s i v t   l � g e   ( e n d a s t   F T P   p r o t o k o l l ) 
     - i m p l i c i t                     I m p l i c i t   T L S / S S L   ( e n d a s t   F T P S   p r o t o k o l l ) 
     - e x p l i c i t s s l               E x p l i c i t   S S L   ( e n d a s t   F T P S   p r o t o k o l l ) 
     - e x p l i c i t t l s               E x p l i c i t   T L S   ( e n d a s t   F T P S   p r o t o k o l l ) 
     - r a w s e t t i n g   s e t t i n g 1 = v � r d e 1   s e t t i n g s 2 = v � r d e 2   . . . 
                                           K o n f i g u r e r a r   v a r j e   s e s s i o n s i n s t � l l n i n g   m e d   r a w - f o r m a t 
                                           s o m   i   e n   I N I - f i l 
 e x e m p e l : 
     o p e n 
     o p e n   s f t p : / / m a r t i n @ e x a m p l e . c o m : 2 2 2 2   - p r i v a t e k e y = m y k e y . p p k 
     o p e n   m a r t i n @ e x a m p l e . c o m 
     o p e n   e x a m p l e . c o m 
 � c l o s e   [   < s e s s i o n >   ] 
     S t � n g e r   s e s s i o n   s p e c i f i c e r a d   m e d   s i t t   n u m m e r .   O m   s e s s i o n s n u m r e t   i n t e   � r 
     s p e c i f i c e r a d ,   s t � n g s   d e n   a k t u e l l a   s e s s i o n e n . 
 e x e m p e l : 
     c l o s e 
     c l o s e   1 
 � s e s s i o n   [   < s e s s i o n >   ] 
     G � r   s e s s i o n e n   s p e c i f i c e r a d   m e d   e t t   n u m m e r   a k t i v .   O m   e t t   s e s s i o n s n u m m e r 
     i n t e   � r   s p e c i f i c e r a d ,   l i s t a s   a n s l u t n a   s e s s i o n e r . 
 e x e m p e l : 
     s e s s i o n 
     s e s s i o n   1 
 ; p w d 
     V i s a r   a k t u e l l   f j � r r k a t a l o g   f � r   d e n   a k t i v a   s e s s i o n e n . 
 � c d   [   < k a t a l o g >   ] 
     � n d r a r   a k t u e l l   k a t a l o g   p �   s e r v e r n   i   d e n   a k t i v a   s e s s i o n e n . 
     O m   e n   k a t a l o g   i n t e   a n g e s ,   a n v � n d s   h e m k a t a l o g e n . 
 e x e m p e l : 
     c d   / h o m e / m a r t i n 
     c d 
 l s   [   < k a t a l o g >   ] / [   < j o k e r t e c k e n > ] 
     V i s a r   i n n e h � l l e t   i   a n g i v e n   f j � r r k a t a l o g .   O m   k a t a l o g   
   i n t e   a n g e s ,   v i s a s   i n n e h � l l e t   i   a k t u e l l   k a t a l o g . 
     N � r   j o k e r t e c k e n   h a r   a n g e t t s ,   t o l k a s   d e t   s o m   e n   g r u p p   f i l e r   s k a   l i s t a s . 
   A n n a r s   l i s t a s   a l l a   f i l e r . 
 a s l i a s : 
     d i r 
 e x e m p e l : 
     l s 
     l s   / h o m e / m a r t i n 
 @ l p w d 
     V i s a r   a k t u e l l   l o k a l   k a t a l o g   ( g � l l e r   f � r   a l l a   s e s s i o n e r ) . 
 J l c d   < k a t a l o g > 
     B y t e r   l o k a l   k a t a l o g   f � r   a l l a   s e s s i o n e r . 
 e x e m p e l : 
     c d   d : \ 
 l l s   [   < k a t a l o g >   ] \ [   < j o k e r t e c k e n >   ] 
     V i s a r   i n n e h � l l e t   i   a n g i v e n   l o k a l   k a t a l o g .   O m   k a t a l o g   
     i n t e   a n g e s ,   v i s a s   i n n e h � l l e t   i   a k t u e l l   k a t a l o g . 
     N � r   j o k e r t e c k e n   h a r   a n g e t t s ,   t o l k a s   d e t   s o m   e n   g r u p p   f i l e r   s k a   l i s t a s . 
   A n n a r s   l i s t a s   a l l a   f i l e r . 
 e x e m p e l : 
     l l s 
     l l s   d : \ 
 r m   < f i l >   [   < f i l 2 >   . . .   ] 
     R a d e r a r   e n   e l l e r   f l e r a   f j � r r f i l e r .   O m   f j � r r p a p p e r s k o r g e n   � r 
     k o n f i g u r e r a d ,   f l y t t a s   f i l e n   d i t   i s t � l l e t   f � r   a t t   r a d e r a s . 
     F i l n a m n   k a n   e r s � t t a s   a v   j o k e r t e c k e n   f � r   a t t   v � l j a   f l e r a   f i l e r . 
 e x e m p e l : 
     r m   i n d e x . h t m l 
     r m   i n d e x . h t m l   a b o u t . h t m l 
     r m   * . h t m l 
 � r m d i r   < k a t a l o g >   [   < k a t a l o g 2 >   . . .   ] 
     R a d e r a r   e n   e l l e r   f l e r a   f j � r r k a t a l o g e r .   O m   f j � r r p a p p e r s k o r g e n   � r 
   k o n f i g u r e r a d ,   f l y t t a s   k a t a l o g e n   d i t   i s t � l l e t   f � r   a t t   r a d e r a s . 
 e x e m p e l : 
     r m d i r   p u b l i c _ h t m l 
  m v   < f i l >   [   < f i l 2 >   . . .   ]   [   < k a t a l o g > /   ] [   < n y t t n a m n >   ] 
     F l y t t a r   e l l e r   b y t e r   n a m n   p �   e n   e l l e r   f l e r a   f j � r r f i l e r .   M � l k a t a l o g e n   e l l e r   n y t t 
     n a m n   e l l e r   b � d a   m � s t e   a n g e s .   M � l k a t a l o g e n   m � s t e   a v s l u t a s   m e d   
     s n e d s t r e c k .   O p e r a t i o n s m a s k   k a n   a n v � n d a s   i s t � l l e t   f � r   n y t t   n a m n . 
     F i l n a m n   k a n   b y t a s   u t   m o t   j o k e r t e c k e n   f � r   a t t   v � l j a   f l e r a   f i l e r . 
 a l i a s : 
     r e n a m e 
 e x e m p e l : 
     m v   i n d e x . h t m l   p u b l c _ h t m l / 
     m v   i n d e x . h t m l   a b o u t . * 
     m v   i n d e x . h t m l   p u b l i c _ h t m l / a b o u t . * 
     m v   p u b l i c _ h t m l / i n d e x . h t m l   p u b l i c _ h t m l / a b o u t . h t m l   / h o m e / m a r t i n / * . b a k 
     m v   * . h t m l   / h o m e / b a c k u p / * . b a k 
 :c h m o d   < m e t o d >   < f i l >   [   < f i l 2 >   . . .   ] 
     � n d r a r   r � t t i g h e t e r n a   p �   e n   e l l e r   f l e r a   f j � r r f i l e r .   M e t o d   k a n   a n g e s 
     s o m   t r e -   e l l e r   f y r s i f f r i g a   o k t a l a   n u m m e r . 
     F i l n a m n   k a n   b y t a s   u t   m o t   j o k e r t e c k e n   f � r   a t t   v � l j a   f l e r a   f i l e r . 
 e x e m p e l : 
     c h m o d   6 4 4   i n d e x . h t m l   a b o u t . h t m l 
     c h m o d   1 7 0 0   / h o m e / m a r t i n / p u b l i c _ h t m l 
     c h m o d   6 4 4   * . h t m l 
 t l n   < m � l >   < s y m b o l i s k   l � n k > 
     S k a p a r   s y m b o l i s k   f j � r r l � n k . 
 a l i a s : 
     s y m l i n k 
 e x e m p e l : 
     l n   / h o m e / m a r t i n / p u b l i c _ h t m l   w w w 
 D m k d i r   < k a t a l o g > 
     S k a p a r   f j � r r k a t a l o g . 
 e x e m p e l : 
     m k d i r   p u b l i c _ h t m l 
 �g e t   < f i l >   [   [   < f i l 2 >   . . .   ]   < k a t a l o g > \ [   < n y t t n a m n >   ]   ] 
     L a d d a r   n e r   e n   e l l e r   f l e r a   f i l e r   f r � n   f j � r r k a t a l o g   t i l l   l o k a l   k a t a l o g . 
     O m   e n d a s t   e n   p a r a m e t e r   a n g e s   l a d d a s   f i l e n   n e r   t i l l   l o k a l 
     a r b e t s k a t a l o g .   O m   f l e r   p a r a m e t r a r   a n g e s ,   a l l a   u t o m   d e n   s i s t a 
     a n g e r   e n   u p p s � t t n i n g   f i l e r   a t t   l a d d a   n e r .   D e n   s i s t a   p a r a m e t e r n   a n g e r   l o k a l 
     m � l k a t a l o g   o c h   e v e n t u e l l   o p e r a t i o n s m a s k   f � r   a t t   s p a r a   f i l e r   u n d e r 
     a n n a t   n a m n .   M � l k a t a l o g e n   m � s t e   s l u t a   m e d   b a c k s l a s h . 
     F i l n a m n   k a n   e r s � t t a s   m e d   j o k e r t e c k e n   f � r   a t t   v � l j a   f l e r a   f i l e r . 
     O m   d u   v i l l   h � m t a   f l e r a   f i l e r   t i l l   a k t u e l l   a r b e t s k a t a l o g   a n v � n d   ' . \ '   s o m 
     s i s t a   p a r a m e t e r n . 
 a l i a s : 
     r e c v ,   m g e t 
 v � x l a r : 
     - d e l e t e                     T a   b o r t   f j � r r k � l l f i l e r   e f t e r   � v e r f � r i n g 
     - r e s u m e                     � t e r u p p t a   � v e r f � r i n g   o m   m � j l i g t   ( e n d a s t   S F T P   o c h   F T P - p r o t o k o l l ) 
     - a p p e n d                     L � g g e r   t i l l   f i l e n   i   s l u t e t   a v   m � l f i l e n   ( e n d a s t   S F T P - p r o t o k o l l ) 
     - p r e s e r v e t i m e         B e v a r a   t i d s s t � m p e l 
     - n o p r e s e r v e t i m e     B e v a r a   i n t e   t i d s s t � m p e l 
     - s p e e d = < k b p s >       B e g r � n s a   � v e r f � r i n g s h a s t i g h e t 
     - t r a n s f e r = < l � g e >   � v e r f � r i n g s l � g e :   b i n a r y ,   a s c i i ,   a u t o m a t i c 
     - f i l e m a s k = < m a s k >   A n g e r   f i l m a s k . 
     - r e s u m e s u p p o r t = < t i l l s t � n d >   K o n f i g u r e r a r   � t e r u p p t a g n i n g s s t � d . 
                                       M � j l i g a   v � r d e n   � r   ' o n ' ,   ' o f f '   e l l e r   t r � s k e l 
 e f f e k t i v a   a l t e r n a t i v : 
     c o n f i r m ,   r e c o n n e c t t i m e 
 e x e m p e l : 
     g e t   i n d e x . h t m l 
     g e t   - d e l e t e   i n d e x . h t m l   a b o u t . h t m l   . \ 
     g e t   i n d e x . h t m l   a b o u t . h t m l   d : \ w w w \ 
     g e t   p u b l i c _ h t m l / i n d e x . h t m l   d : \ w w w \ a b o u t . * 
     g e t   * . h t m l   * . p n g   d : \ w w w \ * . b a k 
 .p u t   < f i l >   [   [   < f i l 2 >   . . .   ]   < k a t a l o g > / [   < n y t t n a m n >   ]   ] 
     � v e r f � r   e n   e l l e r   f l e r a   f i l e r   f r � n   l o k a l   k a t a l o g   t i l l   f j � r r k a t a l o g . 
     O m   e n d a s t   e n   p a r a m e t e r   a n g e s   � v e r f � r s   f i l e n   t i l l   e n   f j � r r a r b e t s k a t a l o g . 
   O m   f l e r a   p a r a m e t r a r   a n g e s ,   a l l a   u t o m   d e n   s i s t a 
     a n g e r   e n   u p p s � t t n i n g   f i l e r   a t t   � v e r f � r a .   D e n   s i s t a   p a r a m e t e r n   a n g e r 
     f j � r r m � l s k a t a l o g   o c h   e v e n t u e l l t   o p e r a t i o n s m a s k   f � r   a t t   s p a r a   f i l e r   u n d e r 
     e t t   a n n a t   n a m n .   M � l k a t a l o g   m � s t e   s l u t a   m e d   e n   s l a s h . 
     F i l n a m n   k a n   e r s � t t a s   m e d   j o k e r t e c k e n   f � r   a t t   v � l j a   f l e r a   f i l e r . 
     F � r   � v e r f � r a   f l e r a   f i l e r   t i l l   a k t u e l l   a r b e t s k a t a l o g ,   a n v � n d   ' . / '   s o m   d e n 
     s i s t a   p a r a m e t e r n . 
 a l i a s : 
     s e n d ,   m p u t 
 v � x l a r : 
     - d e l e t e                           T a   b o r t   l o k a l   k � l l f i l   e f t e r   � v e r f � r i n g 
     - r e s u m e                           � t e r u p p t a   � v e r f � r i n g   o m   m � j l i g t   ( e n d a s t   S F T P   o c h   F T P - p r o t o k o l l ) 
     - a p p e n d                           L � g g   t i l l   f i l   t i l l   s l u t e t   a v   m � l f i l e n   ( e n d a s t   S F T P - p r o t o k o l l ) 
     - p r e s e r v e t i m e               B e v a r a   t i d s s t � m p e l 
     - n o p r e s e r v e t i m e           B e v a r a   i n t e   t i d s s t � m p e l 
     - p e r m i s s i o n s = < l � g e >   A n g e   r � t t i g h e t e r 
     - n o p e r m i s s i o n s             B e h � l l   s t a n d a r d r � t t i g h e t e r 
     - s p e e d = < k i b p s >             B e g r � n s a   � v e r f � r i n g s h a s t i g h e t 
     - t r a n s f e r = < l � g e >         � v e r f � r i n g s l � g e :   b i n a r y ,   a s c i i ,   a u t o m a t i c 
     - f i l e m a s k = < m a s k >         A n g e r   f i l m a s k . 
     - r e s u m e s u p p o r t = < t i l l s t � n d >   K o n f i g u r e r a r   � t e r u p p t a g n i n g s s t � d . 
                                             M � j l i g a   v � r d e n   � r   ' o n ' ,   ' o f f '   e l l e r   t r � s k e l 
 e f f e k t i v a   a l t e r n a t i v : 
     c o n f i r m ,   r e c o n n e c t t i m e 
 e x e m p e l : 
     p u t   i n d e x . h t m l 
     p u t   - d e l e t e   i n d e x . h t m l   a b o u t . h t m l   . / 
     p u t   - p e r m i s s i o n s = 6 4 4   i n d e x . h t m l   a b o u t . h t m l   / h o m e / m a r t i n / p u b l i c _ h t m l / 
     p u t   d : \ w w w \ i n d e x . h t m l   a b o u t . * 
     p u t   * . h t m l   * . p n g   / h o m e / m a r t i n / b a c k u p / * . b a k 
 o p t i o n   [   < a l t e r n a t i v >   [   < v � r d e >   ]   ] 
     O m   i n g a   p a r a m e t r a r   a n g e s ,   v i s a s   a l l a   s c r i p t   a l t e r n a t i v   o c h 
   d e r a s   v � r d e n .   O m   e n d a s t   e n   p a r a m e t e r   a n g e s ,   v i s a s   v � r d e t   f � r   a l t e r n a t i v e t . 
     O m   t v �   p a r a m e t r a r   a n g e s   s � t t   v � r d e t   p �   a l t e r n a t i v e t . 
     U r s p r u n g l i g a   v � r d e n   a v   v i s s a   a l t e r n a t i v   � r   h � m t a d e   f r � n   a p p l i k a t i o n e n s   k o n f i g u r a t i o n , 
     m o d i f i k a t i o n   a v   d e s s a   � n d r a r   d o c k   i n t e   a p p l i k a t i o n e n s 
   k o n f i g u r a t i o n . 
 a l t e r n a t i v   � r : 
     e c h o           o n | o f f 
                       V � x l a r   e k o   a v   k o m m a n d o   s o m   e x e k v e r a s . 
                       P � v e r k a d e   k o m m a n d o n :   a l l 
     b a t c h         o n | o f f | a b o r t | c o n t i n u e 
                       V � x l a r   b a t c h   l � g e   ( a l l a   u p p m a n i n g a r   b e s v a r a s   a u t o m a t i s k t 
                       n e g a t i v t ) .   N � r   ' o n ' ,   r e k o m m e n d e r a s   a t t   s � t t a   ' c o n f i r m ' 
                       t i l l   ' o f f '   f � r   a t t   t i l l � t a   � v e r s k r i v n i n g a r .   M e d   ' a b o r t ' ,   s c r i p t   a v b r y t s 
                       n � r   e t t   f e l   i n t r � f f a r .   M e d   ' c o n t i n u e ' ,   a l l a   f e l   i g n o r e r a s . 
                       P � v e r k a d e   k o m m a n d o n :   n e a r l y   a l l 
     c o n f i r m     o n | o f f 
                       V � x l a r   b e k r � f t e l s e r   ( � v e r s k r i v n i n g ,   e t c . ) . 
                       P � v e r k a d e   k o m m a n d o n :   g e t ,   p u t 
     t r a n s f e r   b i n a r y | a s c i i | a u t o m a t i c 
                       � v e r f � r i n g s l � g e :   b i n a r y ,   a s c i i   ( t e x t ) ,   a u t o m a t i c   ( e f t e r   f i l � n d e l s e ) . 
                       P � v e r k a d e   k o m m a n d o n :   g e t ,   p u t ,   s y n c h r o n i z e ,   k e e p u p t o d a t e 
     e x k l u d e r a     c l e a r   |   < m a s k >   [   ;   < m a s k 2 >   . . .   ] 
     i n k l u d e r a     c l e a r   |   < m a s k >   [   ;   < m a s k 2 >   . . .   ] 
                       S t � l l e r   i n   e x k l u d e r i n g s -   e l l e r   i n k l u d e r i n g s m a s k e r   ( e n d a s t   e n   k a n   v a r a   a k t i v ) . 
                       K a t a l o g e r   p � v e r k a s   o c k s �   ( * /   m a t c h a r   a l l a   k a t a l o g e r ) . 
                       P � v e r k a d e   k o m m a n d o n :   g e t ,   p u t ,   s y n c h r o n i z e ,   k e e p u p t o d a t e 
     r e c o n n e c t t i m e   o f f   |   < s e c > 
                       T i d s b e g r � n s n i n g   i   s e k u n d e r   f � r   � t e r a n s l u t n i n g   a v   b r u t e n   s e s s i o n . 
                       C o m m a n d s   a f f e c t e d :   g e t ,   p u t ,   s y n c h r o n i z e ,   k e e p u p t o d a t e 
 a l i a s e s : 
     a s c i i   =     o p t i o n   t r a n s f e r   a s c i i 
     b i n a r y   =   o p t i o n   t r a n s f e r   b i n a r y 
 e x e m p e l : 
     o p t i o n 
     o p t i o n   t r a n s f e r 
     o p t i o n   c o n f i r m   o f f 
     o p t i o n   i n c l u d e   " * . h t m l ;   * / " 
 As y n c h r o n i z e   l o c a l | r e m o t e | b o t h   [   < l o k a l   k a t a l o g >   [   < f j � r r k a t a l o g >   ]   ] 
     N � r   d e n   f � r s t a   p a r a m e t e r n   � r   ' l o c a l '   s y n k r o n i s e r a s   l o k a l   k a t a l o g   m e d 
     f j � r r k a t a l o g .   N � r   d e n   f � r s t a   p a r a m e t e r n   � r   ' r e m o t e '   s y n k r o n i s e r a s   f j � r r k a t a l o g 
     m e d   l o k a l   k a t a l o g .   N � r   d e n   f � r s t a   p a r a m e t e r n   � r   ' b o t h '   s y n k r o n i s e r a s 
     k a t a l o g e r n a   m o t   v a r a n d r a . 
     N � r   k a t a l o g e r   i n t e   s p e c i f i c e r a s ,   s y n k r o n i s e r a s   a k t u e l l 
     k a t a l o g . 
     O B S :   � v e r s k r i v n i n g s b e k r � f t e l s e r   � r   a l l t i d   a v   f � r   k o m m a n d o t . 
 v � x l a r : 
     - p r e v i e w                           F � r h a n d s g r a n s k a   � n d r i n g a r ,   s y n k r o n i s e r a r   i n t e 
     - d e l e t e                             T a   b o r t   f � r � l d r a d e   f i l e r 
     - m i r r o r                             S p e g e l l � g e   ( s y n k r o n i s e r a r   f � r � l d r a d e   f i l e r   o c k s � ) . 
                                               I g n o r e r a s   m e d   ' b o t h ' . 
     - c r i t e r i a = < k r i t e r i e r >   J � m f � r e l s e k r i t e r i e r .   M � j l i g a   v � r d e n   � r   ' n o n e ' ,   ' t i m e ' , 
                                               ' s i z e '   o c h   ' e i t h e r ' .   I g n o r e r a s   m e d   ' b o t h ' - l � g e . 
     - p e r m i s s i o n s = < l � g e >     A n g e   r � t t i g h e t e r 
     - n o p e r m i s s i o n s               B e h � l l   s t a n d a r d r � t t i g h e t e r 
     - s p e e d = < k b p s >               B e g r � n s a   � v e r f � r i n g s h a s t i g h e t 
     - t r a n s f e r = < l � g e >           � v e r f � r i n g s l � g e :   b i n a r y ,   a s c i i ,   a u t o m a t i c 
     - f i l e m a s k = < m a s k >           A n g e   f i l m a s k . 
     - r e s u m e s u p p o r t = < t i l l s t � n d >   K o n f i g u r e r a r   � t e r u p p t a g n i n g s s t � d . 
                                               M � j l i g a   v � r d e n   � r   ' o n ' ,   ' o f f '   e l l e r   t r � s k e l 
 e f f e k t i v a   a l t e r n a t i v : 
     r e c o n n e c t t i m e 
 e x e m p e l : 
     s y n c h r o n i z e   r e m o t e   - d e l e t e 
     s y n c h r o n i z e   b o t h   d : \ w w w   / h o m e / m a r t i n / p u b l i c _ h t m l 
 ]k e e p u p t o d a t e   [   < l o k a l   k a t a l o g >   [   < f j � r r k a t a l o g >   ]   ] 
     T i t t a r   e f t e r   f � r � n d r i n g a r   i   d e n   l o k a l a   k a t a l o g e n   o c h   � t e r s p e g l a r   d e m   p �   f j � r r k a t a l o g e n . 
     N � r   k a t a l o g e r   i n t e   a n g e s ,   s y n k r o n i s e r a s   a k t u e l l   a r b e t s k a t a l o g 
 .   F � r   a t t   s l u t a   t i t t a   e f t e r   f � r � n d r i n g a r   t r y c k   C t r l - C 
     O B S :   S k r i v a   � v e r   b e k r � f t e l s e r   � r   a l l t i d   a v   f � r   k o m m a n d o t . 
 v � x l a r : 
     - d e l e t e                           T a   b o r t   f � r � l d r a d e   f i l e r 
     - p e r m i s s i o n s = < l � g e >   A n g e   b e h � r i g h e t e r 
     - n o p e r m i s s i o n s             B e h � l l   s t a n d a r d b e h � r i g h e t e r 
     - s p e e d = < k b p s >             B e g r � n s a   � v e r f � r i n g s h a s t i g h e t 
     - t r a n s f e r = < l � g e >         � v e r f � r i n g s l � g e :   b i n a r y ,   a s c i i ,   a u t o m a t i c 
     - f i l e m a s k = < m a s k >         A n g e r   f i l m a s k . 
     - r e s u m e s u p p o r t = < t i l l s t � n d >   K o n f i g u r e r a r   � t e r u p p t a   s t � d . 
                                             M � j l i g a   v � r d e n   � r   ' o n '   o c h   ' o f f '   e l l e r   t r � s k e l 
 e f f e k t i v a   a l t e r n a t i v : 
     r e c o n n e c t t i m e 
 e x e m p e l : 
     k e e p u p t o d a t e   - d e l e t e 
     k e e p u p t o d a t e   d : \ w w w   / h o m e / m a r t i n / p u b l i c _ h t m l 
 Wc a l l   < K o m m a n d o > 
     M e d   S F T P   o c h   S C P   p r o t o k o l l e n ,   k � r s   g o d t y c k l i g t   f j � r r s k a l s k o m m a n d o . 
     O m   a k t u e l l   s e s s i o n   i n t e   t i l l � t e r   k � r n i n g   a v   g o d t y c k l i g   f j � r r k o m m a n d o 
     s k i l d a   s k a l s e s s i o n e r   k o m m e r   a t t   � p p n a s   a u t o m a t i s k t . 
     O m   F T P   p r o t o k o l l ,   k � r   e t t   p r o t o k o l l k o m m a n d o . 
     K o m m a n d o t   k a n   i n t e   k r � v a   a n v � n d a r i n p u t . 
 a l i a s : 
     ! 
 e x e m p e l : 
     c a l l   t o u c h   i n d e x . h t m l 
 ] e c h o   < m e d d e l a n d e > 
     S k r i v e r   m e d d e l a n d e   t i l l   s k r i p t u t d a t a . 
 e x e m p e l : 
     e c h o   S t a r t i n g   u p l o a d . . . 
 Y s t a t   < f i l > 
     H � m t a r   o c h   l i s t a r   a t t r i b u t   f � r   a n g i v e n   f j � r r f i l . 
 e x e m p e l : 
     s t a t   i n d e x . h t m l 
               
 C O R E _ E R R O R " V � r d n y c k e l n   k u n d e   i n t e   v e r i f i e r a s !  A n s l u t n i n g   m i s s l y c k a d e s .  A v s l u t a d   a v   a n v � n d a r e n .  T a p p a d   a n s l u t n i n g . # K a n   i n t e   h i t t a   k o m m a n d o t s   r e t u r k o d . C K o m m a n d o t   ' % s ' 
 m i s s l y c k a d e s   m e d   r e t u r k o d e n   % d   o c h   f e l m e d d e l a n d e 
 % s . ) K o m m a n d o t   m i s s l y c k a d e s   m e d   r e t u r k o d e n   % d . 7 K o m m a n d o t   ' % s '   m i s s l y c k a d e s   m e d   o g i l t i g   u t m a t n i n g   ' % s ' . = F e l   u p p s t o d   n � r   n a m n e t   p �   a k t u e l l   f j � r r k a t a l o g   s k u l l e   h � m t a s . | F e l   u p p s t o d   n � r   s t a r t m e d d e l a n d e   h o p p a d e s   � v e r .   D i t t   s k a l   � r   a n t a g l i g e n   i n k o m p a t i b e l t   m e d   a p p l i k a t i o n e n   ( B A S H   r e k o m m e n d e r a s ) . ) F e l   u p p s t o d   n � r   k a t a l o g   b y t t e s   t i l l   ' % s ' .     ) F e l   u p p s t o d   n � r   l i s t n i n g   a v   k a t a l o g   ' % s ' . % O v � n t a d   k a t a l o g l i s t n i n g   v i d   r a d   ' % s ' . # F e l a k t i g   r � t t i g h e t s b e s k r i v n i n g   ' % s ' ; F e l   u p p s t o d   n � r   d e n   a l l m � n n a   k o n f i g u r a t i o n e n   s k u l l e   r e n s a s . + F e l   u p p s t o d   n � r   l a g r a d e   s e s s i o n e r   r e n s a d e s . 1 F e l   u p p s t o d   n � r   f i l e n   m e d   s l u m p t a l s f r � n   r e n s a d e s . - F e l   u p p s t o d   n � r   c a c h a d e   v � r d n y c k l a r   r e n s a d e s . Q F e l   u p p s t o d   n � r   v a r i a b e l   i n n e h � l l a n d e   r e t u r k o d   a v   s e n a s t e   k o m m a n d o   s k u l l e   h i t t a s . 0 F e l   u p p s t o d   n � r   a n v � n d a r g r u p p e r   s k u l l e   s l � s   u p p . " F i l   e l l e r   k a t a l o g   ' % s '   f i n n s   i n t e . ) K a n   i n t e   h i t t a   a t t r i b u t e n   f � r   f i l e n   ' % s ' .  K a n   i n t e   � p p n a   f i l e n   ' % s ' . ( F e l   u p p s t o d   n � r   f i l e n   ' % s '   s k u l l e   l � s a s . 3 A l l v a r l i g t   f e l   u p p s t o d   v i d   k o p i e r i n g   a v   f i l e n   ' % s ' . 0 F i l k o p i e r i n g e n   t i l l   f j � r r k a t a l o g e n   m i s s l y c k a d e s . 0 F i l k o p i e r i n g e n   f r � n   f j � r r k a t a l o g e n   m i s s l y c k a d e s . % S C P   p r o t o k o l l f e l :   O v � n t a d   r a d b r y t n i n g & S C P   p r o t o k o l l f e l :   F e l a k t i g t   t i d s f o r m a t 2 S C P   p r o t o k o l l f e l :   F e l a k t i g   c o n t r o l   r e c o r d   ( % s ;   % s ) # K o p i e r i n g   a v   f i l   ' % s '   m i s s l y c k a d e s . 1 S C P   p r o t o k o l l f e l :   F e l a k t i g t   f i l b e s k r i v n i n g s f o r m a t  ' % s '   � r   i n g e n   k a t a l o g ! ( F e l   u p p s t o d   n � r   k a t a l o g e n   ' % s '   s k a p a d e s .  K a n   i n t e   s k a p a   f i l e n   ' % s ' . * F e l   u p p s t o d   v i d   s k r i v n i n g   t i l l   f i l e n   ' % s ' . * K a n   i n t e   s � t t a   a t t r i b u t e n   t i l l   f i l e n   ' % s ' . + F e l m e d d e l a n d e   m o t t a g e t   f r � n   f j � r r s i d a :   ' % s ' " F e l   v i d   b o r t t a g n i n g   a v   f i l e n   ' % s ' . 7 F e l   u p p s t o d   v i d   l o g g n i n g   o c h   d e n   h a r   d � r f � r   s t � n g t s   a v .  K a n   i n t e   � p p n a   l o g g f i l e n   ' % s ' . 0 F e l   u p p s t o d   n � r   f i l e n   ' % s '   b y t t e   n a m n   t i l l   ' % s ' .     F i l e n   m e d   n a m n   ' % s '   f i n n s   r e d a n . $ K a t a l o g e n   m e d   n a m n   ' % s '   f i n n s   r e d a n . 2 F e l   u p p s t o d   v i d   b y t e   a v   k a t a l o g   t i l l   h e m k a t a l o g e n . ' F e l   u p p s t o d   v i d   r e n s n i n g   a v   a l l a   a l i a s .   ; F e l   u p p s t o d   n � r   n a t i o n e l l a   a n v � n d a r v a r i a b l e r   s k u l l e   r e n s a s . ! O v � n t a d   i n d a t a   f r � n   s e r v e r n :   ' % s ' ( F e l   u p p s t o d   n � r   I N I - f i l e n   s k u l l e   r e n s a s .   6 A u t e n t i s e r i n g s l o g g   ( s e   s e s s i o n s l o g g   f � r   d e t a l j e r ) : 
 % s 
  A u t e n t i s e r i n g   m i s s l y c k a d e s . # A n s l u t n i n g e n   h a r   o v � n t a t   a v s l u t a t s . 1 F e l   u p p s t o d   n � r   n y c k e l n   s p a r a d e s   t i l l   f i l e n   ' % s ' .   ) S e r v e r n   s k i c k a d e   k o m m a n d o t   s l u t s t a t u s   % d . < S F T P   p r o t o k o l l v a r n i n g :   F e l a k t i g   m e d d e l a n d e t y p   v i d   s v a r   ( % d ) .   I S F T P - s e r v e r n s   v e r s i o n   ( % d )   s t � d s   i n t e .   V e r s i o n e r   s o m   s t � d s   � r   % d   t i l l   % d . E S F T P   p r o t o k o l l v a r n i n g :   F e l a k t i g t   m e d d e l a n d e n u m m e r   % d   ( f � r v � n t a d e   % d ) .  O v � n t a d   O K   r e s p o n s .  O v � n t a d   E O F   r e s p o n s . ! F i l e n   e l l e r   k a t a l o g e n   f i n n s   i n t e .  � t k o m s t   n e k a d . . A l l m � n t   f e l   ( s e r v e r n   b o r d e   g e   f e l b e s k r i v n i n g ) . J D � l i g t   m e d d e l a n d e   ( D � l i g t   f o r m a t e r a t   p a k e t   e l l e r   i n k o m p a t i b e l t   p r o t o k o l l ) .  I n g e n   a n s l u t n i n g .  F � r l o r a d   a n s l u t n i n g .   S e r v e r n   s t � d e r   i n t e   o p e r a t i o n e n . - % s 
 F e l k o d :   % d 
 F e l m e d d e l a n d e   f r � n   s e r v e r % s :   % s  O k � n d   s t a t u s k o d . ' F e l   v i d   l � s n i n g   a v   s y m b o l i s k   l � n k   ' % s ' . 4 S e r v e r n   r e t u r n e r a d e   t o m   l i s t n i n g   f � r   k a t a l o g e n   ' % s ' . 6 M o t t o g   S S H _ F X P _ N A M E   p a k e t   m e d   n o l l   e l l e r   f l e r a   p o s t e r .   + K a n   i n t e   f �   d e n   v e r k l i g a   s � k v � g e n   f � r   ' % s ' . ) K a n   i n t e   � n d r a   e g e n s k a p e r   f � r   f i l e n   ' % s ' . F K a n   i n t e   i n i t i a l i s e r a   S F T P - p r o t o k o l l e t .   K � r   v � r d d a t o r n   e n   S F T P - s e r v e r ? " K a n   i n t e   l � s a   t i d s z o n s i n f o r m a t i o n .  K a n   i n t e   s k a p a   f j � r r f i l   ' % s ' .  K a n   i n t e   � p p n a   f j � r r f i l   ' % s ' .  K a n   i n t e   s t � n g a   f j � r r f i l   ' % s ' .  ' % s '   � r   i n t e   e n   f i l ! � � v e r f � r i n g e n   l y c k a d e s   s l u t f � r a ,   m e n   t e m p o r � r   � v e r f � r i n g s f i l   ' % s '   k u n d e   i n t e   b y t a   n a m n   t i l l   m � l f i l   ' % s ' .   O m   p r o b l e m e t   k v a r s t � r ,   p r o v a   m e d   a t t   s l �   a v   f i l � v e r f � r i n g e n s   � t e r u p p t a - f u n k t i o n  K a n   i n t e   s k a p a   l � n k   ' % s ' .  O g i l t i g t   k o m m a n d o   ' % s ' .  I n g e n 4 ' % s '   � r   i n g e n   t i l l � t e n   f i l r � t t i g h e t   i   o k t a l t   f o r m a t . 5 S e r v e r n   k r � v e r   e t t   e j   s t � t t   s l u t - p � - r a d   s e k v e n s   ( % s ) .  O k � n d   f i l t y p   ( % d )  O g i l t i g t   v e r k t y g .   % S � k v � g e n   f i n n s   i n t e   e l l e r   � r   o g i l t i g .  F i l e n   f i n n s   r e d a n . R F i l e n   l i g g e r   p �   e n   e n h e t   s o m   e n d a s t   s t � d e r   l � s n i n g ,   e l l e r   e n h e t e n   � r   s k r i v s k y d d a d .   D e t   f i n n s   i n g e t   m e d i a   i   e n h e t e n . * F e l   u p p s t o d   v i d   a v k o d n i n g   a v   U T F - 8   s t r � n g . < F e l   u p p s t o d   v i d   k � r n i n g   a v   e g e t   k o m m a n d o   ' % s '   p �   f i l e n   ' % s ' .  K a n   i n t e   l a d d a   l o c a l e   % d . + M o t t o g   e j   k o m p l e t t a   d a t a p a k e t   f � r e   f i l s l u t . 8 F e l   u p p s t o d   v i d   b e r � k n i n g   a v   s t o r l e k   f � r   k a t a l o g e n   ' % s ' . L M o t t o g   e t t   f � r   s t o r t   ( % d   B )   S F T P   p a k e t .   M a x i m a l t   s t � d d   p a k e t s t o r l e k   � r   % d   B . � K a n   i n t e   k � r a   S C P   f � r   a t t   s t a r t a   � v e r f � r i n g .   K o n t r o l l e r a   a t t   S C P   � r   i n s t a l l e r a t   p �   s e r v e r n   o c h   a t t   s � k v � g e n   � r   i n k l u d e r a d   i   P A T H .   D u   k a n   o c k s �   p r o v a   S F T P   i s t � l l e t   f � r   S C P .  P l a t s p r o f i l e n   ' % s '   f i n n s   r e d a n . , F e l   u p p s t o d   v i d   f l y t t   a v   f i l   ' % s '   t i l l   ' % s ' . x % s 
   
 F e l e t   o r s a k a s   n o r m a l t   a v   e t t   m e d d e l a n d e   f r � n   e t t   i n l o g g n i n g s s k r i p t   ( s o m   . p r o f i l e ) .   M e d d e l a n d e t   k a n   s t a r t a   m e d   " % s " . � * * � v e r f � r i n g   a v   f i l   ' % s '   l y c k a d e s ,   m e n   f e l   u p p s t o d   v i d   i n s t � l l n i n g   a v   r � t t i g h e t e r   o c h / e l l e r   t i d s s t � m p e l . * * 
 
 O m   p r o b l e m e t   k v a r s t � r ,   s t � n g   a v   a n g e   r � t t i g h e t e r   e l l e r   b e v a r a   t i d s s t � m p e l .   A l t e r n a t i v e t   k a n   d u   a k t i v e r a   a l t e r n a t i v e t   ' I g n o r e r a   r � t t i g h e t s f e l ' .  O g i l t i g   � t k o m s t   t i l l   m i n n e t .   2 D e t   f i n n s   i n g e n   l e d i g t   u t r y m m e   k v a r   i   f i l s y s t e m e t . t O p e r a t i o n e n   k a n   i n t e   s l u t f � r a s   p �   g r u n d   a v   a t t   d e t   s k u l l e   m e d f � r a   a t t   a n v � n d a r e n s   l a g r i n g s - q u o t a   s k u l l e   � v e r s k r i d a s . $ P r i n c i p a l   ( % s )   � r   o k � n t   f � r   s e r v e r n . 0 F e l   u p p s t o d   v i d   k o p i e r i n g   a v   f i l   ' % s '   t i l l   ' % s ' . ( O a v s l u t a t   m � n s t e r   ' % s '   v i d   b � r j a n   a v   % d . $ O k � n t   m � n s t e r   ' % s '   v i d   b � r j a n   a v   % d . V K a n   i n t e   k o m b i n e r a   f i l n a m n s m � n s t e r   ( b � r j a r   v i d   % d )   m e d   f i l l i s t m � n s t e r   ( b � r j a r   v i d   % d ) .  O k � n t   k o m m a n d o   ' % s ' . 0 T v e t y d i g t   k o m m a n d o   ' % s ' .   M � j l i g   m a t c h n i n g   � r :   % s $ P a r a m e t e r   s a k n a s   f � r   k o m m a n d o t   ' % s ' . ( F � r   m � n g a   p a r a m e t r a r   f � r   k o m m a n d o t   ' % s ' .          I n g e n   s e s s i o n .  O g i l t i g t   s e s s i o n s n u m m e r   ' % s ' .  O k � n t   a l t e r n a t i v   ' % s ' . % O k � n t   v � r d e   ' % s '   f � r   a l t e r n a t i v   ' % s ' . ( K a n   i n t e   b e s t � m m a   s t a t u s   p �   s o c k e t   ( % d ) . � F e l   u p p s t o d   v i d   b o r t t a g n i n g   a v   f i l   ' % s ' .   E f t e r   � t e r u p p t a g e n   f i l � v e r f � r i n g   m � s t e   b e f i n t l i g   m � l f i l   t a s   b o r t .   O m   d u   i n t e   h a   r � t t i g h e t e r   a t t   t a   b o r t   m � l f i l ,   m � s t e   d u   a v a k t i v e r a   � t e r u p p t a g n i n g   a v   f i l � v e r f � r i n g . 5 F e l   u p p s t o d   v i d   a v k o d n i n g   a v   S F T P   p a k e t   ( % d ,   % d ,   % d ) . 1 O g i l t i g t   n a m n   ' % s ' .   N a m n   k a n   i n t e   i n n e h � l l a   ' % s ' . @ F i l e n   k u n d e   i n t e   � p p n a s   f � r   a t t   d e n   � r   l � s t   a v   e n   a n n a n   p r o c e s s .  K a t a l o g e n   � r   i n t e   t o m . + D e n   s p e c i f i c e r a d e   f i l e n   � r   i n t e   e n   k a t a l o g .  F i l n a m n e t   � r   i n t e   g i l t i g t . ( F � r   m � n g a   s y m b o l i s k a   l � n k a r   a n t r � f f a d e s .  F i l e n   k a n   i n t e   t a s   b o r t . p E n   a v   p a r a m e t r a r n a   v a r   u t a n f � r   i n t e r v a l l e t ,   e l l e r   p a r a m e t r a r n a   s o m   s p e c i f i c e r a d e s   k a n   i n t e   a n v � n d a s   t i l l s a m m a n s . V D e n   s p e c i f i c e r a d e   f i l e n   v a r   e n   k a t a l o g ,   i   e n   k o n t e x t   d � r   e n   k a t a l o g   i n t e   k a n   a n v � n d a s .  L � s   f � r   b y t e i n t e r v a l l   k r o c k a d e .    L � s   f � r   b y t e i n t e r v a l l   n e k a d e s . P E n   o p e r a t i o n   f � r s � k t e   g � r a s   p �   e n   f i l   s o m   h a r   e n   v � n t a n d e   b o r t t a g n i n g s o p e r a t i o n . F F i l e n   � r   k o r r u p t ;   e n   k o n t r o l l   a v   i n t e g r i t e t e n   i   f i l s y s t e m e t   b � r   k � r a s . L F i l e n   ' % s '   f i n n s   i n t e   e l l e r   d e n   i n n e h � l l e r   i n t e   p r i v a t   n y c k e l   i   k � n t   f o r m a t . � P r i v a t   n y c k e l f i l   ' % s '   i n n e h � l l e r   n y c k e l   i   % s   f o r m a t .   W i n S C P   s t � d e r   b a r a   P u T T Y   f o r m a t . 
   
 D u   k a n   a n v � n d a   P u T T Y g e n   v e r k t y g e t   f � r   a t t   k o n v e r t e r a   d i n   p r i v a t a   n y c k e l f i l . i P r i v a t   n y c k e l f i l   ' % s '   i n n e h � l l e r   n y c k e l   i   % s   f o r m a t .   D e n   f � l j e r   i n t e   d i n   f � r e d r a g n a   S S H   p r o t o k o l l v e r s i o n . { K a n   i n t e   s k r i v a   � v e r   f j � r r f i l   ' % s ' . 
   
 T r y c k   ' T a   b o r t '   f � r   a t t   t a   b o r t   f i l   o c h   s k a p a   e n   n y   i s t � l l e t   f � r   a t t   s k r i v a   � v e r   d e n .  & T a   b o r t = F e l   u p p s t o d   v i d   k o n t r o l l   a v   l e d i g t   u t r y m m e   f � r   s � k v � g e n   ' % s ' . S K a n   i n t e   h i t t a   l e d i g   l o k a l   l i s t n i n g s p o r t n u m m e r   f � r   t u n n e l   i   i n t e r v a l l e t   % d   t i l l   % d . * K a n   i n t e   u t f � r a   n � t v e r k s h � n d e l s e   ( f e l   % d ) . / S e r v e r n   a v s l u t a d e   o v � n t a t   n � t v e r k s a n s l u t n i n g e n . 1 F e l   u p p s t o d   n � r   a n s l u t n i n g e n   s k u l l e   t u n n l a s . 
   
 % s 9 F e l   u p p s t o d   n � r   k o n t r o l l s u m m a n   b e r � k n a d e s   f � r   f i l e n   ' % s ' .  I n t e r n t   f e l   % s   ( % s ) .  O p e r a t i o n e n   s t � d s   i n t e .    � t k o m s t   n e k a d . ' F r � g a r   e f t e r   a u t e n t i s e r i n g s u p p g i f t e r . . . $ O g i l t i g   s v a r   t i l l   P W D   k o m m a n d o   ' % s ' . + T h i s   v e r s i o n   d o e s   n o t   s u p p o r t   F T P   p r o t o c o l .  O k � n d   v � x e l   ' % s ' . ) F e l   u p p s t o d   v i d   � v e r f � r i n g   a v   f i l e n   ' % s ' .  K a n   i n t e   k � r a   ' % s ' .  F i l e n   ' % s '   h i t t a d e s   i n t e . . E t t   f e l   u p p s t o d   n � r   d o k u m e n t e t   s k u l l e   s t � n g a s . % ' % s '   � r   i n g e n   g i l t i g   h a s t i g h e t s g r � n s .  C e r t i f i c a t e   c h a i n   t o o   l o n g .  C e r t i f i c a t e   h a s   e x p i r e d .  C e r t i f i c a t e   i s   n o t   y e t   v a l i d .  C e r t i f i c a t e   r e j e c t e d .  C e r t i f i c a t e   s i g n a t u r e   f a i l u r e .  C e r t i f i c a t e   n o t   t r u s t e d .  S j � l v s i g n e r a t   c e r t i f i k a t . , F o r m a t   f e l   i   c e r t i f i k a t e t s   g i l t i g - t i l l   f � l t . , F o r m a t   f e l   i   c e r t i f i k a t e t s   g i l t i g - f r � n   f � l t .  O g i l t i g   C A   c e r t i f i k a t .  E j   s t � t t   c e r t i f i k a t   � n d a m � l . 5 N y c k e l a n v � n d n i n g   i n k l u d e r a r   i n t e   c e r t i f i k a t s i g n e r i n g . , B e g r � n s n i n g a r   f � r   s � k v � g s l � n g d e n   � v e r s k r i d s . + S j � l v s i g n e r a t   c e r t i f i k a t   i   c e r t i f i k a t k e d j a . 6 D e t   g � r   i n t e   a t t   a v k o d a   u t f � r d a r e n s   o f f e n t l i g a   n y c k e l . 3 D e t   g � r   i n t e   a t t   d e k r y p t e r a   c e r t i f i k a t e t s   s i g n a t u r . + D e t   g � r   i n t e   a t t   f �   u t f � r d a r e n s   c e r t i f i k a t . 2 D e t   g � r   i n t e   a t t   h � m t a   l o k a l t   u t f � r d a t   c e r t i f i k a t . 3 D e t   g � r   i n t e   a t t   v e r i f i e r a   d e t   f � r s t a   c e r t i f i k a t e t . % O k � n t   f e l   v i d   k o n t r o l l   a v   c e r t i f i k a t . 6 F e l e t   i n t r � f f a d e   p �   e t t   d j u p   a v   % d   i   c e r t i f i k a t k e d j a n .      M a s k e n   � r   o g i l t i g   n � r a   ' % s ' . � S e r v e r n   k a n   i n t e   � p p n a   a n s l u t n i n g   i   a k t i v t   l � g e .   O m   d u   s i t t e r   b a k o m   e n   N A T - r o u t e r ,   k a n   d u   b e h � v a   a n g e   e n   e x t e r n   I P - a d r e s s .   A l t e r n a t i v t ,   � v e r v � g a   a t t   b y t a   t i l l   p a s s i v t   l � g e . ( F e l   u p p s t o d   v i d   b o r t t a g n i n g   a v   f i l   ' % s ' . ? O g i l t i g t   v � r d e   p �   v � x e l   ' % s ' .   G i l t i g a   v � r d e n   � r   ' o n '   o c h   ' o f f ' .  � t k o m s t   u t a n   l � s e n o r d   n e k a d . 0 K a n   i n t e   � p p n a   w e b b p l a t s k a t a l o g   e l l e r   a r b e t s y t a . ) N � t v e r k s f e l :   I n g e   v � g   t i l l   v � r d   " % H O S T % " . 2 N � t v e r k s f e l :   M j u k v a r a   o r s a k a d e   a v b r u t e n   a n s l u t n i n g  V � r d   " % H O S T % "   f i n n s   i n t e . 0 I n k o m m a n d e   p a k e t   v a r   f � r v a n s k a t   v i d   d e k r y p t e r i n g U % s 
 
 H j � l p   o s s   a t t   f � r b � t t r a   W i n S C P   g e n o m   a t t   r a p p o r t e r a   f e l   p �   W i n S C P : s   s u p p o r t f o r u m . - F e l   v i d   a v k o d n i n g   a v   T L S / S S L - c e r t i f i k a t   ( % s ) .  C O R E _ C O N F I R M A T I O N M V � r d e n   k o m m u n i c e r a r   i n t e   u n d e r   % d   s e k u n d e r . 
 
 V � n t a   y t t e r l i g a r e   % 0 : d   s e k u n d e r ?    & L � s e n o r d   f � r   n y c k e l n   ' % s ' : # F i l e n   ' % s '   f i n n s   r e d a n .   S k r i v   � v e r ? ' K a t a l o g e n   ' % s '   f i n n s   r e d a n .   S k r i v   � v e r ? � D e t   f � r s t a   % s s k i f f r e t   s o m   s t � d s   a v   s e r v e r n   � r   % s ,   s o m   l i g g e r   u n d e r   k o n f i g u r e r a d   v a r n i n g s t r � s k e l n . 
 
 V i l l   d u   f o r t s � t t a   m e d   d e n   h � r   a n s l u t n i n g e n ?    k l i e n t - t i l l - s e r v e r  s e r v e r - t i l l - k l i e n t � * * V i l l   d u   � t e r u p p t a   f i l � v e r f � r i n g e n ? * * 
 
 M � l k a t a l o g e n   i n n e h � l l e r   d e l v i s   � v e r f � r d   f i l   ' % s ' . 
 
 O B S : S v a r a   ' N e j '   t a r   b o r t   d e l v i s   � v e r f � r d   f i l   o c h   s t a r t a r   o m   � v e r f � r i n g . o M � l k a t a l o g e n   i n n e h � l l e r   d e n   d e l v i s   � v e r f � r d a   f i l e n   ' % s ' ,   s o m   � r   s t � r r e   � n   k � l l f i l e n .   F i l e n   k o m m e r   a t t   t a s   b o r t . u * * V i l l   d u   l � g g a   t i l l   f i l e n   ' % s '   i   s l u t e t   a v   b e f i n t l i g   f i l ? * * 
 
 T r y c k   ' N e j '   f � r   a t t   � t e r u p p t a   f i l � v e r f � r i n g e n   i s t � l l e t . 4 % s 
   
 N y :             	 % s   b y t e s ,   % s 
 B e f i n t l i g :   	 % s   b y t e s ,   % s ' F i l e n   ' % s '   � r   s k r i v s k y d d a d .   S k r i v   � v e r ? � * * S k r i v   � v e r   l o k a l   f i l   ' % s ' ? * * M � l k a t a l o g e n   i n n e h � l l e r   r e d a n   f i l e n   ' % s ' . 
 V � l j   o m   d u   v i l l   s k r i v a   � v e r   f i l e n   e l l e r   h o p p a   � v e r   d e n n a   � v e r f � r i n g   o c h   b e h � l l a   b e f i n t l i g   f i l . � * * S k r i v   � v e r   f j � r r f i l   ' % s ' ? * * M � l k a t a l o g e n   i n n e h � l l e r   r e d a n   f i l e n   ' % s ' . 
 V � l j   o m   d u   v i l l   s k r i v a   � v e r   f i l e n   e l l e r   h o p p a   � v e r   d e n n a   � v e r f � r i n g   o c h   b e h � l l a   b e f i n t l i g   f i l .         � V � r d   k o m m u n i c e r a r   i n t e   m e r   � n   n � g r a   ' % d '   s e k u n d e r .   V � n t a r   f o r t f a r a n d e . . . 
 
 O B S :   O m   p r o b l e m e t   u p p r e p a s ,   p r o v a   a t t   s t � n g a   a v   ' O p t i m e r a   s t o r l e k e n   p �   a n s l u t n i n g s b u f f e r t ' . � D e n   f � r s t a   a l g o r i t m e n   f � r   n y c k e l u t b y t e   s o m   s t � d s   a v   s e r v e r n   � r   % s ,   s o m   l i g g e r   u n d e r   k o n f i g u r e r a d   v a r n i n g s t r � s k e l . 
 
 V i l l   d u   f o r t s � t t a   m e d   d e n   h � r   a n s l u t n i n g e n ?  & � t e r a n s l u t 
 N y t t   n a & m n      T u n n e l   f � r   % s  L � s e n o r d  L � s e n o r d   f � r   n y c k e l  S e r v e r p r o m p t  A n v � n d a r n a m n  A & n v � n d a r n a m n :  S e r v e r p r o m p t :   % s  N y t t   l � s e n o r d  S & v a r :    A n v � n d e r   T I S   a u t e n t i s e r i n g . % s $ A n v � n d e r   K r y p t o k o r t   a u t e n t i s e r i n g . % s 
 & L � s e n o r d : / A n v � n d e r   t a g e n t b o r d s i n t e r a k t i v   a u t e n t i s e r i n g . % s  N & u v a r a n d e   l � s e n o r d :  & N y t t   l � s e n o r d  & B e k r � f t a   n y t t   l � s e n o r d :  A u t e n t i s e r i n g   f � r   t u n n e l s e s s i o n  � v e r f � r   m e d   e t t   a n n a t   n a m n  & N y t t   n a m n : g* * S e r v e r n s   c e r t i f i k a t   � r   i n t e   k � n t .   D u   h a r   i n g e n   g a r a n t i   f � r   a t t   s e r v e r n   � r   d e n   d a t o r   s o m   d u   t r o r   a t t   d e   � r . * * 
 
 S e r v e r c e r t i f i k a t e t s   d e t a l j e r   f � l j e r : 
 
 % s 
 
 O m   d u   l i t a r   p �   c e r t i f i k a t e t ,   t r y c k   p �   ' J a ' .   F � r   a t t   a n s l u t a   u t a n   a t t   l a g r a   c e r t i f i k a t   t r y c k e r   d u   p �   ' N e j ' .   F � r   a t t   a v b r y t a   a n s l u t n i n g e n   t r y c k e r   p �   A v b r y t . 
 
 V i l l   d u   f o r t s � t t a   a n s l u t a   o c h   l a g r a   c e r t i f i k a t e t ? - -   O r g a n i s a t i o n :   % s 
 | -   P l a t s :   % s 
 | -   A n n a t :   % s 
  % s ,   % s S U t g i v a r e : 
 % s 
 � m n e : 
 % s 
 G i l t i g :   % s   -   % s 
 
 F i n g e r a v t r y c k   ( S H A 1 ) :   % s 
 
 S a m m a n f a t t n i n g :   % s                        F i l n a m n   f � r   c e r t i f i k a t  A n g e   f i l n a m n   f � r   c e r t i f i k a t :              C O R E _ I N F O R M A T I O N  J a  N e j G V � r d :   % s 
 A n v � n d a r n a m n :   % s 
 P r i v a t   n y c k e l f i l :   % s 
 � v e r f � r i n g s p r o t o k o l l :   % s  V e r s i o n   % d . % d . % d   ( B y g g d   % d ) > O p e r a t i o n e n   s l u t f � r d e s   f r a m g � n g s r i k t .   A n s l u t n i n g e n   a v s l u t a d e s .  S F T P - % d : S F T P   p r o t o k o l l e t s   v e r s i o n   t i l l � t e r   i n t e   n a m n b y t e   p �   f i l e r . ' S e r v e r n   s t � d e r   i n g a   u t � k n i n g a r   a v   S F T P . ( S e r v e r n   s t � d e r   f � l j a n d e   S F T P   u t � k n i n g a r :     
 L � & g g   t i l l  E n d a s t   n & y a r e  V i s a r   h j � l p . S t � n g e r   a l l a   s e s s i o n e r   o c h   a v s l u t a r   p r o g r a m m e t    A n s l u t e r   t i l l   s e r v e r  S t � n g e r   s e s s i o n e n 4 L i s t a r   a n s l u t n a   s e s s i o n e r   e l l e r   v � l j e r   a k t i v   s e s s i o n  V i s a r   a k t u e l l   f j � r r k a t a l o g  B y t e r   a k t u e l l   f j � r r k a t a l o g  V i s a r   i n n e h � l l e t   i   f j � r r k a t a l o g  V i s a r   a k t u e l l   l o k a l   k a t a l o g  B y t e r   a k t u e l l   l o k a l   k a t a l o g ! L i s t a r   i n n e h � l l e t   i   l o k a l   k a t a l o g  T a r   b o r t   f j � r r f i l  T a r   b o r t   f j � r r k a t a l o g $ F l y t t a r   e l l e r   b y t e r   n a m n   p �   f j � r r f i l   � n d r a r   r � t t i g h e t e r n a   p �   f j � r r f i l  S k a p a r   e n   s y m b o l i s k   f j � r r l � n k  S k a p a r   f j � r r k a t a l o g 3 L a d d a r   n e r   f i l   f r � n   f j � r r k a t a l o g   t i l l   l o k a l   k a t a l o g 3 L a d d a r   u p p   f i l   f r � n   l o k a l   k a t a l o g   t i l l   f j � r r k a t a l o g - S � t t e r   e l l e r   v i s a r   v � r d e n   p �   s c r i p t a l t e r n a t i v , S y n k r o n i s e r a r   f j � r r k a t a l o g   m e d   l o k a l   k a t a l o g D K o n t i n u e r l i g t   � t e r s p e g l a   � n d r i n g a r   i   l o k a l   k a t a l o g   t i l l   f j � r r k a t a l o g  V � r d :      A k t i v   s e s s i o n :   [ % d ]   % s  S e s s i o n   ' % s '   a v s l u t a d .  L o k a l   ' % s '   % s   F j � r r   ' % s '  ' % s '   b o r t t a g e n 7 � v e r v a k a r   f � r � n d r i n g a r ,   t r y c k   C T R L - C   f � r   a t t   a v b r y t a . . .  & H o p p a   � v e r   a l l a  K � r   g o d t y c k l i g t   f j � r r k o m m a n d o  & T e x t  & B i n � r t   8 � v e r f � r i n g s t y p :   % s | B i n � r | T e x t | A u t o m a t i s k   ( % s ) | A u t o m a t i s k O F i l n a m n s f � r � n d r i n g :   % s | I n g e n   � n d r i n g | V e r s a l e r | G e m e n e r | F � r s t a   v e r s a l | G e m e n e r   8 . 3  S � t t   r � t t i g h e t e r :   % s  L � g g   t i l l   X   t i l l   k a t a l o g  B e v a r a   t i d s s t � m p e l    F i l m a s k :   % s  R e n s a   ' A r k i v '   a t t r i b u t  B y t   i n t e   u t   o g i l t i g a   t e c k e n    B e v a r a   i n t e   t i d s s t � m p e l  B e r � k n a   i n t e   � v e r f � r i n g s s t o r l e k   S t a n d a r d � v e r f � r i n g s i n s t � l l n i n g a r  V � r d n a m n :   % s  A n v � n d a r n a m n :   % s  F j � r r k a t a l o g :   % s    L o k a l   k a t a l o g :   % s $ S k a n n a r   ' % s '   e f t e r   u n d e r k a t a l o g e r . . . % � v e r v a k a r   � n d r i n g a r   i   % d   k a t a l o g e r . . .  � n d r i n g   i   ' % s '   u p p t � c k t .  F i l   ' % s '   � v e r f � r d .  F i l   ' % s '   b o r t t a g e n . U % s   k o n f i g u r e r a d   � v e r f � r i n g s i n s t � l l n i n g   k a n   i n t e   a n v � n d a s   i   a k t u e l l   k o n t e x t | N � g o n | A l l a    I g n o r e r a   r � t t i g h e t s f e l  A n v � n d e r   a n v � n d a r n a m n   " % s " . . A n v � n d e r   t a n g e n t b o r d s i n t e r a k t i v   a u t e n t i s e r i n g . % A u t e n t i s e r i n g   m e d   p u b l i k   n y c k e l   " % s " .  F e l a k t i g   l � s e n o r d .  � t k o m s t   n e k a d . 0 A u t e n t i s e r i n g   m e d   p u b l i k   n y c k e l   " % s "   f r � n   a g e n t . ( F � r s � k e r   m e d   p u b l i k   n y c k e l a u t e n t i s e r i n g . ' A u t e n t i s e r i n g   m e d   f � r i n s t � l l t   l � s e n o r d .  � p p n a r   t u n n e l . . .  A n s l u t n i n g   a v s l u t a d .    S � k e r   e f t e r   v � r d . . .  A n s l u t e r   t i l l   v � r d . . .  A u t e n t i s e r a r . . .  A u t e n t i s e r a d .  S t a r t a r   s e s s i o n e n . . .  L � s e r   f j � r r k a t a l o g . . .  S e s s i o n e n   s t a r t a d .  A n s l u t e r   g e n o m   t u n n e l . . .  S e r v e r   n e k a r   v � r   n y c k e l .  A d m i n i s t r a t i v t   f � r b j u d e n   ( % s ) .  A n s l u t n i n g   m i s s l y c k a d e s   ( % s ) . . N � t v e r k s f e l :   A n s l u t n i n g   t i l l   " % H O S T % "   n e k a d e s .   + N � t v e r k s f e l :   A n s l u t n i n g   � t e r s t � l l d   a v   p e e r . 5 N � t v e r k s f e l :   A n s l u t n i n g   t i l l   " % H O S T % "   g j o r d e   t i m e o u t . 2 V � r d :   % s 
 A n v � n d a r n a m n :   % s 
 � v e r f � r i n g s p r o t o k o l l :   % s 
 & � t e r u p p t a / S e r v e r n   s t � d e r   i n t e   n � g r a   e x t r a   F T P   e g e n s k a p e r . . S e r v e r n   s t � d e r   d e   h � r   e x t r a   F T P   e g e n s k a p e r n a :   # � v e r f � r i n g s h a s t i g h e t s g r � n s :   % u   k B / s  & K o p i e r a   n y c k e l 
 & U p p d a t e r a 
 & L � g g   t i l l  B e v a r a   e n d a s t   l � s n i n g 	 J � m f � r . . .  S y n k r o n i s e r a r . . .  I n g e t   a t t   s y n k r o n i s e r a . 
 O b e g r � n s a d  S S L / T L S   I m p l i c i t   k r y p t e r i n g    S S L   E x p l i c i t   k r y p t e r i n g  T L S   E x p l i c i t   k r y p t e r i n g  V i s a r   a r g u m e n t e n   s o m   m e d d e l a n d e  H � m t a r   a t t r i b u t   f � r   f j � r r f i l # V � r d e n s   f i n g e r a v t r y c k s n y c k e l   � r   % s . F V � x e l   - f i l e m a s k   � s i d o s � t t e r   f � r � l d r a d e   i n k l u d e r a / e x k l u d e r a   a l t e r n a t i v .  B a r a   & n y a   o c h   � n d r a d e   f i l e r � S e r v e r n   a v v i s a d e   S F T P - a n s l u t n i n g ,   m e n   d e n   l y s s n a r   p �   F T P - a n s l u t n i n g a r . 
 
 V i l l   d u   a n v � n d a   F T P - p r o t o k o l l e t   i s t � l l e t   f � r   S F T P ?   F � r e d r a r   a t t   a n v � n d a   k r y p t e r i n g . ` � p p n a   s e s s i o n   m e d   k o m m a n d o r a d s p a r a m e t e r   i   s k r i p t   � r   f � r � l d r a d .   A n v � n d   ' o p e n ' - k o m m a n d o t   i s t � l l e t . L V A R N I N G !   A t t   g e   u p p   s � k e r h e t e n   o c h   a c c e p t e r a   n � g o n   n y c k e l   s o m   k o n f i g u r e r a t s ! P V A R N I N G !   A t t   g e   u p p   s � k e r h e t e n   o c h   a c c e p t e r a   n � g o t   c e r t i f i k a t   s o m   k o n f i g u r e r a t s !  N y   l o k a l   f i l   % s  N y   f j � r r f i l   % s $ L o k a l   f i l   % s   � r   n y a r e   � r   f j � r r f i l   % s $ F j � r r f i l   % s   � r   n y a r e   � n   l o k a l   f i l   % s  � v e r g e   f j � r r f i l   % s    � v e r g e   l o k a l   f i l   % s  S k i l l n a d e r   h i t t a d e :  T a   b o r t   E O F - t e c k e n  T a   b o r t   B O M                                            C O R E _ V A R I A B L E ( S S H   o c h   S C P   k o d e n   � r   b a s e r a d   p �   P u T T Y   % s  0 . 6 3 " C o p y r i g h t   �   1 9 9 7 - 2 0 1 3   S i m o n   T a t h a m 2 h t t p : / / w w w . c h i a r k . g r e e n e n d . o r g . u k / ~ s g t a t h a m / p u t t y /  F T P - k o d   b a s e r a d   p �   F i l e Z i l l a    C o p y r i g h t   �   T i m   K o s s e  h t t p : / / f i l e z i l l a - p r o j e c t . o r g / m D e n n a   p r o d u k t   i n n e h � l l e r   p r o g r a m v a r a   s o m   u t v e c k l a t s   a v   O p e n S S L   P r o j e c t   f � r   a n v � n d n i n g   i   O p e n S S L : s   v e r k t y g   % s . ) C o p y r i g h t   �   1 9 9 8 - 2 0 1 4   T h e   O p e n S S L   P r o j e c t  1 . 0 . 1 h  h t t p : / / w w w . o p e n s s l . o r g /                         > h t t p : / / w w w . c h i a r k . g r e e n e n d . o r g . u k / ~ s g t a t h a m / p u t t y / l i c e n c e . h t m l            * *                                         $ E r r o r   r e t r i e v i n g   f i l e   l i s t   f o r   " % s " . n C e r t i f i c a t e   w a s   n o t   i s s u e d   f o r   t h i s   s e r v e r .   Y o u   m i g h t   b e   c o n n e c t i n g   t o   a   s e r v e r   t h a t   i s   p r e t e n d i n g   t o   b e   " % s " .                         �D u   f � r s � k e r   f l y t t a   f j � r r f i l e r   t i l l   e n   d e s t i n a t i o n   s o m   W i n S C P   i n t e   d i r e k t   k a n   f l y t t a   t i l l .   F i l e r n a   k o m m e r   a t t   l a d d a s   n e r   t i l l   e n   t e m p o r � r   k a t a l o g   i s t � l l e t .   A n s v a r e t   f � r   � v e r f � r i n g e n   t i l l   d e n   s l u t g i l t i g a   d e s t i n a t i o n e n   s k a   s k � t a s   a v   m � l a p p l i k a t i o n e n   ( t .   e x .   U t f o r s k a r e n ) ,   v i l k e t   W i n S C P   i n t e   k a n   k o n t r o l l e r a .   K � l l f i l e r   k o m m e r   a t t   r a d e r a s   e f t e r   a t t   n e r l a d d n i n g e n   t i l l   d e n   t e m p o r � r a   k a t a l o g e n   h a r   a v s l u t a t s .   O m   m � l a p p l i k a t i o n e n   m i s s l y c k a s   m e d   a t t   h a n t e r a   d e   t e m p o r � r a   f i l e r n a ,   k a n   d e   f � r l o r a s .   � v e r v � g   g � r n a   a t t   k o p i e r a   f i l e r n a   i s t � l l e t   f � r   a t t   f l y t t a   d e m . 
 T i p s :   F � r   a t t   k o p i e r a   f i l e r   h � l l   n e r   C T R L   t a n g e n t e n   m e d a n   f l y t t . 
 
 V i l l   d u   f o r t f a r a n d e   f l y t t a   f i l e r n a ? [W i n S C P ,   % s 
 % s 
 
 A n v � n d n i n g : 
 G : % A P P %   s e s s i o n 
 G : % A P P %   [ ( s f t p | s c p | f t p ) : / / ] [ a n v � n d a r e [ : l � s e n o r d ] @ ] v � r d [ : p o r t ] [ / s � k v � g / [ f i l ] ] 
 G : % A P P %   [ s e s s i o n ]   / s y n c h r o n i z e   [ l o k a l _ d i r ]   [ f j � r r _ d i r ]   [ / d e f a u l t s ] 
 G : % A P P %   [ s e s s i o n ]   / k e e p u p t o d a t e   [ l o k a l _ d i r ]   [ f j � r r _ d i r ]   [ / d e f a u l t s ] 
 G : % A P P %   [ s e s s i o n ]   / p r i v a t e k e y = < n y c k e l >   / h o s t k e y = < f i n g e r a v t r y c k > 
 G : % A P P %   [ s e s s i o n ]   / c e r t i f i c a t e = < f i n g e r a v t r y c k >   / i m p l i c i t | e x p l i c i t s s l | e x p l i c i t t l s 
 G : % A P P %   [ s e s s i o n ]   / p a s s i v e = o n | o f f   / t i m e o u t = < s e k > 
 G : % A P P %   [ s e s s i o n ]   / r a w s e t t i n g s   s e t t i n g 1 = v � r d e 1   s e t t i n g s 2 = v � r d e 2   . . . 
 G : % A P P %   [ / c o n s o l e ]   [ / s c r i p t = f i l ]   [ / c o m m a n d   k o m m a n d o 1 . . . ]   [ / p a r a m e t e r   p a r a m e t e r 1 . . . ] 
 C : % A P P %   [ / s c r i p t = f i l ]   [ / c o m m a n d   k o m m a n d o 1 . . . ]   [ / p a r a m e t e r   p a r a m e t e r 1 . . . ] 
 B : % A P P %   / i n i = < i n i - f i l >   / l o g = < l o g g f i l >   / x m l l o g = < l o g g f i l > 
 G : % A P P %   / u p d a t e 
 B : % A P P %   / h e l p 
 
 G :   s e s s i o n               N a m n   p �   s p a r a d   s e s s i o n   e l l e r   d i r e k t   s e s s i o n - s p e c i f i k a t i o n . 
 G :   / s y n c h r o n i z e     S y n k r o n i s e r a r   i n n e h � l l e t   i   t v �   k a t a l o g e r . 
 G :   / k e e p u p t o d a t e   S t a r t s   H � l l e r   f j � r r k a t a l o g   a k t u e l l   f u n k t i o n . 
 G :   / d e f a u l t s           S t a r t a r   o p e r a t i o n   u t a n   a t t   v i s a   d i a l o g r u t a . 
 G :   / c o n s o l e             K o n s o l l � g e   ( t e x t ) .   S t a n d a r d l � g e ,   n � r   d e t   a n r o p a s 
 G :                               a n v � n d e r   % A P P % . c o m . 
 B :   / s c r i p t =             K � r   k o m m a n d o f i l .   O m   s k r i p t e t   i n t e   s l u t a r   m e d 
 B :                               ' e x i t '   k o m m a n d o ,   n o r m a l t   i n t e r a k t i v t   l � g e   f � l j e r . 
 B :   / c o m m a n d             K � r   l i s t a   m e d   s k r i p t k o m m a n d o n . 
 B :   / p a r a m e t e r         S k i c k a r   l i s t a   m e d   p a r a m e t r a r   t i l l   s k r i p t . 
 B :   / i n i =                   S � k v � g   t i l l   k o n f i g u r a t i o n   I N I - f i l . 
 B :   / l o g =                   S � t t e r   p �   s e s s i o n s l o g g n i n g   t i l l   f i l . 
 B :   / x m l l o g =             S � t t e r   p �   X M L - l o g g n i n g   t i l l   f i l . 
 G :   / p r i v a t e k e y =     P r i v a t   n y c k e l f i l . 
 G :   / t i m e o u t =           S e r v e r s v a r e t s   t i m e o u t . 
 G :   / h o s t k e y =           F i n g e r a v t r y c k   f � r   s e r v e r n s   v � r d n y c k e l . 
 G :   / p a s s i v e =           P a s s i v t   l � g e   ( e n d a s t   F T P   p r o t o k o l l ) . 
 G :   / r a w s e t t i n g s =   K o n f i g u r e r a r   v a r j e   s e s s i o n s i n s t � l l n i n g   m e d   r a w - f o r m a t 
 G :                               s o m   i   e n   I N I - f i l . 
 G :   / c e r t i f i c a t e =   F i n g g e r a v t r y c k   f � r   S S L / T L S   c e r t i f i k a t . 
 G :   / i m p l i c i t           I m p l i c i t   T L S / S S L   ( e n d a s t   F T P S   p r o t o k o l l ) . 
 G :   / e x p l i c i t s s l     E x p l i c i t   S S L   ( e n d a s t   F T P S   p r o t o k o l l ) . 
 G :   / e x p l i c i t t l s     E x p l i c i t   T L S   ( e n d a s t   F T P S   p r o t o k o l l ) . 
 G :   / u p d a t e               F r � g a r   a p p l i k a t i o n e n s   h e m s i d a n   o m   u p p d a t e r i n g a r . 
 B :   / h e l p                   S k r i v e r   d e t t a   m e d d e l a n d e . 
                                   	 W I N _ E R R O R   Q % s 
   
 V a r n i n g :   A t t   a v b r y t a   d e n   h � r   o p e r a t i o n e n   k o m m e r   a t t   s t � n g a   n e r   a n s l u t n i n g e n !          K a n   i n t e   s k a p a   g e n v � g . ) K a n   i n t e   s k r i v a   � v e r   s p e c i a l s e s s i o n   ' % s ' .  K a n   i n t e   u t f o r s k a   k a t a l o g   ' % s ' . + I n g e n   f i l l i s t a   f � r   � v e r f � r i n g   h a r   a n g i v i t s .  K a n   i n t e   s k a p a   k a t a l o g e n   ' % s ' .   ' K a n   i n t e   t a   b o r t   t e m p o r � r   k a t a l o g   ' % s ' . % K a n   i n t e   � p p n a   e l l e r   k � r a   f i l e n   ' % s ' .  K a n   i n t e   s t a r t a   e d i t o r   ' % s ' .   w K a n   i n t e   � p p n a   m o t s v a r a d e   k a t a l o g   i   m o t s a t t   p a n e l .   S y n k r o n i s e r i n g   a v   k a t a l o g b l � d d r i n g   m i s s l y c k a d e s .   D e n   h a r   s t � n g t s   a v .  K a n   i n t e   a v g � r a   g e n v � g   ' % s ' .   % ' % s '   � r   i n t e   g i l t i g t   p r o f i l p l a t s n a m n . 4 ' % s '   � r   i n t e   g i l t i g t   n a m n   f � r   e n   p r o f i l p l a t s k a t a l o g . 1 P r o f i l p l a t s k a t a l o g e n   m e d   n a m n e t   ' % s '   f i n n s   r e d a n . 5 B e s k r i v n i n g   p �   e g e t   k o m m a n d o   k a n   i n t e   i n n e h � l l a   ' % s ' . 1 E g e t   k o m m a n d o   m e d   b e s k r i v n i n g e n   ' % s '   f i n n s   r e d a n . D K a n   i n t e   f r � g a   a p p l i k a t i o n e n s   h e m s i d a   e f t e r   u p p d a t e r i n g s i n f o r m a t i o n . , F e l   u p p s t o d   v i d   s � k n i n g   e f t e r   u p p d a t e r i n g a r .         < K a n   i n t e   r e g i s t r e r a   p r o g r a m m e t   f � r   a t t   h a n t e r a   U R L - a d r e s s e r . 2 M u t e x   s l � p p t e s   i n t e   e n l i g t   d e t   k r � v d a   i n t e r v a l l e t . E S k a l   d r a - t i l l � g g e t   m u t e x   s l � p p t e s   i n t e   e n l i g t   d e t   k r � v d a   i n t e r v a l l e t . �* * W i n S C P   k u n d e   i n t e   i d e n t i f i e r a   k a t a l o g e n ,   s o m   f i l e n   s l � p p t e s   i . * *   A n t i n g e n   h a r   d u   i n t e   s l � p p t   f i l e n   i   e n   v a n l i g   k a t a l o g   ( t . e x .   U t f o r s k a r e n )   e l l e r   o m   d u   i n t e   h a r   s t a r t a t   o m   d a t o r n   � n n u   e f t e r   i n s t a l l a t i o n e n   a v   s k a l t i l l � g g e t   d r a   &   s l � p p . 
 
 A l t e r n a t i v t   k a n   d u   v � x l a   t i l l   k o m p a t i b e l   d r a   &   s l � p p l � g e   ( f r � n   i n s t � l l n i n g s f � n s t r e t ) ,   s o m   a n v � n d e r   t e m p o r � r a   k a t a l o g e r   f � r   n e d l a d d n i n g a r .   D e t   g � r   a t t   d u   s l � p p a   f i l e r   t i l l   a l l a   d e s t i n a t i o n e r . K F i l e n   ' % s '   i n n e h � l l e r   i n t e   n � g o n   � v e r s � t t n i n g   f � r   d e n   h � r   p r o d u k t v e r s i o n e n .   5 F i l e n   ' % s '   i n n e h � l l e r   � v e r s � t t n i n g   f � r   % s   v e r s i o n   % s . � * * D r a   &   s l � p p   s k a l t i l l � g g e t   � r   a k t i v t ,   m e n   t i l l � g g e t   � r   i n t e   i n s t a l l e r a t . * *   I n s t a l l e r a   t i l l � g g e t   e l l e r   b y t   t i l l   k o m p a t i b e l   d r a   &   s l � p p l � g e   ( f r � n   i n s t � l l n i n g s f � n s t r e t ) ,   s o m   a n v � n d e r   t e m p o r � r a   k a t a l o g e r   f � r   n e d l a d d n i n g . 8 G S S A P I / S S P I   m e d   K e r b e r o s   s t � d s   i n t e   p �   d e t   h � r   s y s t e m e t . ' F e l   u p p s t o d   v i d   b e v a k n i n g   a v   � n d r i n g a r . 8 F e l   u p p s t o d   v i d   b e v a k n i n g   a v   � n d r i n g a r   i   k a t a l o g e n   ' % s ' .   6 F e l   u p p s t o d   v i d   b e v a k n i n g e n   a v   � n d r i n g a r   i   f i l e n   ' % s ' . � * * K a n   i n t e   � v e r f � r a   d e n   r e d i g e r a d e   f i l e n   ' % s ' * * 
 
 S e s s i o n e n   ' % s '   h a r   r e d a n   s t � n g t s . 
 
 � p p n a   e n   n y   s e s s i o n   p �   s a m m a   w e b b p l a t s   o c h   f � r s � k   s p a r a   f i l e n   i g e n . I D e t   f i n n s   r e d a n   f � r   m � n g a   f i l e r   � p p n a d e .   V a r   g o d   s t � n g   n � g r a   f i l e r   f � r s t .   R % s   V a r   v � n l i g   t a   b o r t   f i l e n .   A n n a r s   k o m m e r   i n t e   a p p l i k a t i o n e n   a t t   f u n g e r a   k o r r e k t . o K a n   i n t e   s k a p a   t e m p o r � r   k a t a l o g   ' % s ' .   D u   k a n   � n d r a   r o t k a t a l o g e n   f � r   l a g r i n g   a v   t e m p o r � r a   f i l e r   i   I n s t � l l n i n g a r . �W i n S C P   k u n d e   i n t e   a v g � r a   v i l k e t   p r o g r a m   s o m   s k a   s t a r t a s   f � r   a t t   � p p n a   f i l e n .   W i n S C P   k a n   i n t e   b e v a k a   � n d r i n g a r   i   f i l e n ,   s �   d e n   v i l l   i n t e   l a d d a s   u p p . 
   
 E n   m � j l i g   o r s a k   t i l l   p r o b l e m e t   � r   a t t   f i l e n   r e d a n   h a r   � p p n a t s   a v   e t t   a n n a t   p r o g r a m   s o m   k � r s . 
   
 O m   d u   v i l l   a n v � n d a   p r o g r a m m e t   f � r   a t t   � p p n a   f i l e r   f r � n   W i n S C P ,   � v e r v � g   a t t   k o n f i g u r e r a   d e n   s o m   e n   e x t e r n   e d i t o r . 
   
 N o t e r a   a t t   f i l e n   l i g g e r   k v a r   i   d e n   t e m p o r � r a   k a t a l o g e n . � N � g r a   a v   d e   t e m p o r � r a   k a t a l o g e r n a   k u n d e   i n t e   t a s   b o r t .   O m   f i l e r   f i n n s   l a g r a d e   d � r   s o m   f o r t f a r a n d e   � r   � p p n a ,   s t � n g   d e s s a   o c h   p r o v a   i g e n . � F � r   a t t   a n v � n d a   v a l t   e g e t   k o m m a n d o ,   f � r   b a r a   e n   f i l   v a r a   m a r k e r a d   i   d e n   e n a   p a n e l e n ,   f � r   a t t   k � r a   k o m m a n d o t   p �   d e   v a l d a   f i l e r n a   i   m o t s a t t   p a n e l .   A l t e r n a t i v t   k a n   s a m m a   a n t a l   f i l e r   m a r k e r a s   i   b � d a   p a n e l e r n a   f � r   a t t   k � r a   k o m m a n d o t   p �   m a t c h a n d e   p a r   a v   f i l e r . W F � r   a t t   a n v � n d a   v a l t   e g e t   k o m m a n d o t   f � r   b a r a   e n   f i l   v a r a   m a r k e r a d   i   d e n   l o k a l a   p a n e l e n .   � N � g r a   a v   d e   v a l d a   f j � r r f i l e r n a   l a d d a d e s   i n t e   n e r .   D e t   v a l d a   e g n a   k o m m a n d o t   m � s t e   k � r a s   p �   m a t c h a n d e   p a r   a v   f i l e r ,   v i l k e t   d � r f � r   i n t e   � r   m � j l i g t . $ K a n   i n t e   i n i t i a l i s e r a   e x t e r n   k o n s o l .   N K a n   i n t e   � p p n a   m a p p n i n g s o b j e k t   f � r   a t t   s t a r t a   k o m m u n i k a t i o n   m e d   e x t e r n   k o n s o l . ; T i m e o u t   v � n t a r   p �   e x t e r n   k o n s o l   f � r   a t t   s l u t f � r a   k o m m a n d o t . 4 I n k o m p a t i b e l t   p r o t o k o l l v e r s i o n   f � r   e x t e r n   k o n s o l   % d . D F e l   u p p s t o d   n � r   s � k v � g   ' % s '   l a d e s   t i l l   m i l j � v a r i a b e l   p a t h ( % % P A T H % % ) . H F e l   u p p s t o d   n � r   s � k v � g   ' % s '   t o g s   b o r t   f r � n   m i l j � v a r i a b e l   p a t h ( % % P A T H % % ) .   [ F i l e n   ' % s '   � r   r e d a n   � p p n a d   i   e n   e x t e r n   e d i t o r   ( a p p l i k a t i o n )   e l l e r   h � l l e r   p �   a t t   l a d d a s   u p p . 8 D u   h a r   i n t e   a n g i v i t   n � g o n   a u t o m a t i s k t   v a l   a v   m a s k r e g l e r . D F � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g   m e d   b e s k r i v n i n g   ' % s '   f i n n s   r e d a n . K E g e t   k o m m a n d o   ' % s '   k a n   i n t e   k � r a s   j u s t   n u .   V � l j   f � r s t   f i l e r   t i l l   k o m m a n d o t . A K a n   i n t e   l a d d a   o m   f i l e n   ' % s ' ,   s e s s i o n e n   ' % s '   h a r   r e d a n   a v s l u t a t s .   S A u t o m a t i s k a   � t g � r d e r   � r   a v s t � n g d a   n � r   U R L   a d r e s s e n   t i l l h a n d a h � l l s   p �   k o m m a n d o r a d e n .     L � s e n o r d e t   k a n   i n t e   d e k r y p t e r a s . 3 D u   h a r   i n t e   a n g e t t   k o r r e k t   n u v a r a n d e   h u v u d l � s e n o r d . 0 N y a   o c h   u p p r e p a d e   h u v u d l � s e n o r d e t   � r   i n t e   s a m m a .   F E x t e r n   k o n s o l u t d a t a   d i r i g e r a s   t i l l   p i p e .   S e   t i l l   a t t   p i p e n   l � s e s   f r � n . ) ' % s '   � r   a r b e t s y t a ,   i n t e   w e b b p l a t s k a t a l o g . ) ' % s '   � r   w e b b p l a t s k a t a l o g ,   i n t e   a r b e t s y t a . ) F e l   v i d   e x e k v e r i n g   a v   k o m m a n d o   " % s "   ( % s ) . A K a n   i n t e   l � g g a   t i l l   s � k v � g   t i l l   % P A T H % ,   % P A T H %   � r   r e d a n   f � r   l � n g .                          W I N _ C O N F I R M A T I O N . S e s s i o n   m e d   n a m n   ' % s '   f i n n s   r e d a n .   S k r i v   � v e r ? ! K a t a l o g e n   ' % s '   f i n n s   i n t e .   S k a p a ?  * * A v b r y t   a k t u e l l   � t g � r d ? * * � * * A v b r y t   f i l � v e r f � r i n g ? 
 
 O p e r a t i o n e n   k a n   i n t e   a v b r y t a s   i   m i t t e n   a v   f i l � v e r f � r i n g . 
 T r y c k   ' J a '   f � r   a t t   a v b r y t a   f i l � v e r f � r i n g   o c h   s t � n g a   a n s l u t n i n g e n . 
 T r y c k   ' N e j '   F � r   a t t   a v s l u t a   a k t u e l l   f i l � v e r f � r i n g . 
 T r y c k   ' A v b r y t '   f � r   a t t   f o r t s � t t a   o p e r a t i o n e n . . � r   d u   s � k e r   p �   a t t   d u   v i l l   t a   b o r t   f i l e n   ' % s ' ? 7 � r   d u   s � k e r   p �   a t t   d u   v i l l   t a   b o r t   d e   % d   v a l d a   f i l e r n a ? / A v s l u t a   s e s s i o n e n   ' % s '   o c h   s t � n g   a p p l i k a t i o n e n ?  F r � g a   m i & g   a l d r i g   i g e n 9F � r   l i t e   l e d i g t   u t r y m m e   p �   t e m p o r � r   e n h e t ! 
 
 N � r   f i l e r   d r a s   f r � n   e n   f j � r r k a t a l o g ,   l a d d a s   f i l e r n a   f � r s t   n e r   t i l l   e n   t e m p o r � r   k a t a l o g   ' % s ' .   D e t   � r   % s   l e d i g t   p �   e n h e t e n .   T o t a l   s t o r l e k   f � r   d e   v a l d a   f i l e r n a   � r   % s . 
 
 O B S :   T e m p o r � r   k a t a l o g e n   k a n   � n d r a s   i   I n s t � l l n i n g s f � n s t r e t . 
 
 V i l l   d u   f o r t s � t t a   m e d   a t t   l a d d a   n e r   f i l e r n a ?   ( L � g g   t i l l   k a t a l o g e n   ' % s '   t i l l   b o k m � r k e n ?   - S k a p a   g e n v � g   p �   s k r i v b o r d e t   f � r   s e s s i o n   ' % s ' ? 2 A n v � n d   a k t u e l l a   s e s s i o n s i n t � l l n i n g a r   s o m   s t a n d a r d ?  & H o p p a   � v e r # F i l e n   h a r   � n d r a t s .   S p a r a   � n d r i n g a r ? 9 S k a p a   u t f o r s k a r e n s   ' S k i c k a   t i l l ' - g e n v � g   f � r   s e s s i o n   ' % s ' ?  S k a p a   v a l d   i k o n / g e n v � g ? / A v s l u t a   a l l a   s e s s i o n e r   o c h   s t � n g   a p p l i k a t i o n e n ?   T a   b o r t   v a l d   p r o f i l p l a t s k a t a l o g ?  & F � r e g � e n d e  & N � s t a   3 V i l l   d u   r e g i s t r e r a   W i n S C P   a t t   h a n t e r a   U R L - a d r e s s e r ? L V i l l   d u   r e n s a   u p p   d a t a   f r � n   d e n   h � r   d a t o r n   s o m   h a r   s k a p a t s   a v   a p p l i k a t i o n e n ? ! % s 
 
 V i l l   d u   s t � n g a   a p p l i k a t i o n e n ? G % % s 
 
 V i l l   d u   a v s l u t a   % d   � t e r s t � e n d e   s e s s i o n e r   o c h   s t � n g a   a p p l i k a t i o n e n ? � * * D e t   f i n n s   f o r t f a r a n d e   n � g r a   � v e r f � r i n g a r   i   b a k g r u n d s k � n .   V i l l   d u   k o p p l a   n e r   i a l l a f a l l ? * * 
 
 V a r n i n g :   O m   d u   t r y c k e r   p �   ' O K '   k o m m e r   a l l a   � v e r f � r i n g a r   a t t   a v s l u t a s   o m e d e l b a r t . * * V i l l   d u   � p p n a   s e p a r a t   s k a l s e s s i o n ? * * 
 
 N u v a r a n d e   s e s s i o n   % s   s t � d e r   i n t e   k o m m a n d o t   d u   b e g � r .   S e p a r a t   s k a l s e s s i o n   k a n   � p p n a s   f � r   a t t   b e a r b e t a   k o m m a n d o t . 
 
 O B S :   S e r v e r n   m � s t e   e r b j u d a   U n i x - l i k n a n d e   s k a l   o c h   s k a l e t   m � s t e   a n v � n d a   s a m m a   s � k v � g s s y n t a x   s o m   n u v a r a n d e   s e s s i o n   % s . � D e t   f i n n s   n � g r a   � p p n a   f i l e r .   V a r   v � n l i g   s t � n g   d e m   i n n a n   a p p l i k a t i o n e n   a v s l u t a s . 
   
 O B S :   O m   d e t t a   i n t e   u t f � r s ,   k a n   r e d i g e r a d e   f i l e r   l i g g a   k v a r   i   d e n   t e m p o r � r a   k a t a l o g e n . '* * V i l l   d u   t a   b o r t   t i d i g a r e   t i l l f � l l i g a   k a t a l o g e r ? * * 
 
 W i n S C P   h a r   h i t t a t   % d   t e m p o r � r a   k a t a l o g e r ,   s o m   f � r m o d l i g e n   h a r   s k a p a t s   t i d i g a r e .   D e s s a   k a t a l o g e r   k a n   i n n e h � l l a   f i l e r   s o m   t i d i g a r e   h a r   r e d i g e r a t s   e l l e r   l a d d a t s   n e r . 
 
 D u   k a n   o c k s �   � p p n a   k a t a l o g e r   f � r   a t t   s e   � v e r   i n n e h � l l e t   o c h   t a   b o r t   d e m   s j � l v .  & � p p n a # V i s a   i n t e   d e t   h � r   m e d d e l a n d e t   i & g e n   f * * V i l l   d u   s k a p a   s k r i v b o r d s i k o n   f � r   a l l a   a n v � n d a r e ? * * 
 
 D u   m � s t e   h a   a d m i n i s t r a t � r s r � t t i g h e t e r   f � r   d e t t a . U V i l l   d u   l � g g a   t i l l   a p p l i k a t i o n e n s   s � k v � g   ' % s '   t i l l   m i l j � v a r i a b e l n s   s � k v � g   ( % % P A T H % % ) ? �E d i t o r n   ( a p p l i k a t i o n )   s o m   s t a r t a d e s   f � r   a t t   � p p n a   f i l   ' % s '   a v s l u t a d e s   f � r   t i d i g t .   O m   d e n   i n t e   a v s l u t a d e s   a v   e r ,   k a n   d e t   b e r o   p �   a t t   d e n   e x t e r n a   e d i t o r   � p p n a r   f l e r a   f i l e r   i   e t t   f � n s t e r   ( p r o c e s s ) .   Y t t e r l i g a r e   s t a r t a d e   i n s t a n s e r   a v   e d i t o r n   s k i c k a r   s e d a n   d e n   n y a   f i l e n   t i l l   b e f i n t l i g a   i n s t a n s e r   a v   e d i t o r n   o c h   a v s l u t a r   s i g   o m e d e l b a r t .   F � r   a t t   s t � d j a   d e n n a   t y p   a v   e d i t o r s ,   m � s t e   W i n S C P   a n p a s s a   s i t t   b e t e e n d e ,   i n t e   t a   b o r t   t e m p o r � r   f i l   n � r   p r o c e s s e n   a v s l u t a r ,   u t a n   a t t   b e h � l l a   d e n   s �   l � n g e   W i n S C P   � r   i g � n g .   B e t e e n d e t   k a n   s t � n g a s   a v   g e n o m   a t t   � n d r a   i n s t � l l n i n g a r   f � r   e d i t o r n   ' E x t e r n   e d i t o r   � p p n a r   v a r j e   f i l   i   e t t   s e p a r a t   f � n s t e r   ( p r o c e s s ) ' .   O m   d i n   e d i t o r   i n t e   � r   a v   d e t   h � r   s l a g e t ,   b o r t s e   f r � n   d e t t a   m e d d e l a n d e   o c h   l � t   f i l e n   t a s   b o r t   f r � n   d e n   t e m p o r � r a   k a t a l o g e n   n u . 
   
 V i l l   n i   t a   b o r t   d e n   � p p n a d e   f i l e n   n u ?   ( G e n o m   a t t   t r y c k a   p �   ' N e j '   k o m m e r   d u   a t t   m � j l i g g � r a   d e t   s � r s k i l d a   b e t e e n d e t   o c h   b e h � l l a   f i l e n   i   t e m p o r � r a   k a t a l o g e n . )   � * * V i l l   d u   g � r a   r i k t n i n g e n   d u   v a l t   t i l l   s t a n d a r d ? * * 
 
 D u   h a r   � s i d o s a t t   f � r v a l d   s y n k r o n i s e r i n g s r i k t n i n g .   S o m   s t a n d a r d   b e s t � m s   r i k t n i n g e n   a v   f i l p a n e l e n   s o m   v a r   a k t i v   i n n a n   i n n a n   d u   k � r d e   s y n k r o n i s e r i n g s f u n k t i o n e n . � * * V i l l   d u   f � r s t   u t f � r a   e n   f u l l s t � n d i g   s y n k r o n i s e r i n g   a v   f j � r r k a t a l o g e n ? * * 
 
 F u n k t i o n e n   ' H � l l   f j � r r k a t a l o g   u p p d a t e r a d '   f u n g e r a r   k o r r e k t   e n d a s t   o m   f j � r r k a t a l o g e n   � r   s y n k r o n i s e r a d   m e d   d e n   l o k a l a   i n n a n   d e n   s t a r t a r . 1 S � k e r   p �   a t t   d u   v i l l   t a   b o r t   s p a r a d   s e s s i o n   ' % s ' ? � F l e r   � n   % d   k a t a l o g e r   o c h   u n d e r k a t a l o g e r   h i t t a d e s .   B e v a k n i n g   a v   � n d r i n g a r   i   m � n g a   k a t a l o g e r   k a n   s i g n i f i k a n t   m i n s k a   p r e s t a n d a n   p �   d a t o r n . 
   
 V i l l   d u   s k a n n a   f l e r   k a t a l o g e r ,   u p p   t i l l   % d   k a t a l o g e r ? 	 % s   ( % d   s )   8 S � k e r   p �   a t t   d u   v i l l   f l y t t a   f i l   ' % s '   t i l l   p a p p e r s k o r g e n ? > S � k e r   p �   a t t   d u   v i l l   f l y t t a   % d   v a l d a   f i l e r   t i l l   p a p p e r s k o r g e n ? I F i l e n   h a r   � n d r a t s .   � n d r i n g a r   v i l l   f � r l o r a s ,   o m   f i l e n   l a d d a s   o m .   F o r t s � t t ?  K & o n f i g u r e r a . . . ^ * * V i l l   d u   f � r s � k a   s k a p a   k a t a l o g e n   ' % s ' ? * * 
 
 K a n   i n t e   � p p n a   m o t s v a r a n d e   k a t a l o g   i   m o t s a t t   p a n e l .  L � g g   t i l l   & d e l a d e   b o k m � r k e n s* * V i l l   d u   s k i c k a   m e d d e l a n d e t   t i l l   W i n S C P : s   w e b b p l a t s ? * * 
 
 D e t   f i n n s   i n g e n   h j � l p s i d a   a s s o c i e r a d   m e d   m e d d e l a n d e t .   W i n S C P   k a n   s � k a   p �   s i n   d o k u m e n t a t i o n s p l a t s   e f t e r   m e d d e l a n d e t e x t e n . 
 
 O B S :   W i n S C P   k o m m e r   a t t   s k i c k a   m e d d e l a n d e t   � v e r   e n   o s � k e r   a n s l u t n i n g .   K o n t r o l l e r a   a t t   m e d d e l a n d e t   i n t e   i n n e h � l l e r   n � g o n   d a t a   s o m   d u   v i l l   s k y d d a ,   t i l l   e x e m p e l   n a m n   p �   f i l e r ,   k o n t o n   e l l e r   v � r d a r . 9* * D i t t   l � s e n o r d   � r   f � r   e n k e l t   o c h   k a n   i n t e   g e   t i l l r � c k l i g t   s k y d d   m o t   a t t a c k e r   m e d   o r d l i s t a   e l l e r   b r u t e   f o r c e . 
 � r   d u   s � k e r   a t t   d u   v i l l   a n v � n d a   d e t ? * * 
 
 O B S :   b r a   l � s e n o r d   h a r   m i n s t   s e x   t e c k e n   o c h   i n n e h � l l e r   b � d e   g e m e n e r   o c h   v e r s a l e r ,   s i f f r o r   o c h   s p e c i a l t e c k e n ,   s �   s o m   a v g r � n s a r e ,   s y m b o l e r ,   b o k s t � v e r   m e d   a c c e n t ,   e t c . 9 S k a p a   g e n v � g   p �   s k r i v b o r d e t   t i l l   w e b b p l a t s k a t a l o g e n   ' % s ' ? 0 S k a p a   g e n v � g   p �   s k r i v b o r d e t   t i l l   a r b e t s y t a   ' % s ' ? E V i l l   d u   � t e r a n s l u t a   s e s s i o n   ' % s '   f � r   a t t   � v e r f � r a   r e d i g e r a d   f i l   ' % s ' ? � * * A v s l u t a   a l l a   s e s s i o n e r   o c h   s t � n g   p r o g r a m m e t   u t a n   a t t   s p a r a   a r b e t s y t a ? * * 
 
 T r y c k   ' N e j '   f � r   a t t   a k t i v e r a   a u t o m a t i s k   s p a r a n d e   a v   a r b e t s y t a . l A n p a s s a d   t e x t r e d i g e r a r e   ' % s '   u p p t � c k t e s . 
 
 V i l l   d u   a n v � n d a   ' % s '   i s t � l l e t   f � r   d e n   i n t e r n a   s t a n d a r d r e d i g e r a r e n ? � * * D u   h a r   s p a r a t   s e s s i o n e r / w e b b p l a t s e r   i   % s . 
 
 V i l l   d u   i m p o r t e r a   d e m   t i l l   W i n S C P ? * * 
 
 ( D u   k a n   i m p o r t e r a   d e m   n � r   s o m   h e l s t   s e n a r e   i   d i a l o g r u t a n   L o g g a   i n ) | P u T T Y   S S h - k l i e n t | F i l e z i l l a   F T P - k l i e n t | % s   o c h   % s k I m p o r t e r a   k o n f i g u r a t i o n   k o m m e r   a t t   s k r i v a   � v e r   a l l a   d i n a   i n s t � l l n i n g a r   o c h   w e b b p l a t s e r . 
 
 V i l l   d u   f o r t s � t t a ?  & A l l a    J & a   t i l l   a l l a  R a & p p o r t e r a � D e t   f i n n s   a n d r a   i n s t a n s e r   a v   W i n S C P   i g � n g . 
 
 S t � l l a   i n   e l l e r   r e n s a   h u v u d l � s e n o r d e t ,   m e d a n   e n   a n n a n   i n s t a n s   a v   W i n S C P   � r   i g � n g ,   k a n   o r s a k a   f � r l u s t   a v   d i n a   l a g r a d e   l � s e n o r d . 
 
 V � n l i g e n   a v s l u t a   a n d r a   i n s t a n s e r   a v   W i n S C P   i n n a n   d u   f o r t s � t t e r . � V i l l   d u   b i f o g a   r e d i g e r a d   f i l   ' % s '   t i l l   s e s s i o n   ' % s ' ? * * 
 
 O r i g i n a l   s e s s i o n e n   s o m   a n v � n d e s   f � r   a t t   l a d d a   n e r   f i l e n   ' % s '   t i l l   e d i t o r n   h a r   r e d a n   s t � n g t s . @ V i l l   d u   a v r e g i s t r e r a   W i n S C P   f r � n   h a n t e r i n g   a v   a l l a   U R L - a d r e s s e r ?                                          W I N _ I N F O R M A T I O N  % s   -   % s  I n g a   s k i l l n a d e r   h i t t a d e s .  � p p n a r   s e s s i o n   ' % s ' 
 % s ' V � n t a r   p �   a t t   d o k u m e n t e t   s k a   s t � n g a s . . .  % s   ( � v e r f � r   m e d   S F T P   e l l e r   S C P )  % s   ( � v e r f � r   m e d   S F T P   e l l e r   S C P )  L o k a l :   % s 
 F j � r r :   % s    & T o u c h  & K � r     1 % d   f e l   u p p s t o d   v i d   s e n a s t e   o p e r a t i o n e n .   V i s a   d e m ?  F e l   % d   a v   % d : 
 % s  D u   h a r   d e n   s e n a s t e   v e r s i o n e n .  N y   v e r s i o n   % s   h a r   s l � p p t s . ! ' % s '   v � r d e   p �   k o m m a n d o & p a r a m e t e r :  ' % s '   k o m m a n d o p a r a m e t e r                        U R L :   P r o t o k o l l e t   % s  A n s l u t e r . . .  F r � g a  F e l  P r o m p t 	 V � n t a r . . .  T a & r / G Z i p . . .  & A r k i v n a m n :  & U n T a r / G Z i p . . .  P a c k a   & u p p   t i l l   k a t a l o g :  & J � m f � r   f i l e r  & G r e p . . .    & S � k   e f t e r   m � n s t e r :  % d   L � s e r   k a t a l o g  B e r � k n a r . . .  
   
 % s 
 L a d d a   & n e r  & K o n t r o l l e r a   i g e n ; F � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g   ' % s '   v a l d e s   a u t o m a t i s k t . 4 � t e r g �   t i l l   f � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g   ' % s ' . + � t e r g �   t i l l   s t a n d a r d � v e r f � r i n g s i n s t � l l n i n g .  R e g e l   f � r   a u t o m a t i s k t   v a l : 
 % s    A d   H o c  P a u s a  & I n t e r n   e d i t o r �A p p l i k a t i o n   s t a r t a d   f � r   a t t   � p p n a   f i l   ' % s '   s t � n g d e s   f � r   t i d i g t .   O m   d e n   i n t e   s t � n g d e s   a v   d i g ,   d e   k a n   b e r o   p �   a t t   a p p l i k a t i o n e n   � p p n a r   f l e r a   f i l e r   i   e t t   f � n s t e r   ( p r o c e s s ) .   Y t t e r l i g a r e   s t a r t a d e   i n s t a n s e r   a v   a p p l i k a t i o n e n   s k i c k a r   d �   d e n   n y a   f i l e n   t i l l   b e f i n t l i g   a p p l i k a t i o n   o c h   s t � n g s   o m e d e l b a r t .   W i n S C P   k a n   s t � d j a   s � d a n a   a p p l i k a t i o n e r   e n d a s t   s o m   e x t e r n   e d i t o r . 
   
 O m   d u   v i l l   a n v � n d a   a p p l i k a t i o n e n   f � r   a t t   � p p n a   f i l e r   f r � n   W i n S C P ,   � v e r v � g a   a t t   k o n f i g u r e r a   d e n   s o m   e n   e x t e r n   e d i t o r .   = R e d i g e r a   ( e x t e r n ) | R e d i g e r a   v a l d a   f i l e r   m e d   e x t e r n   e d i t o r   ' % s ' � *   m a t c h a r   a l l a   a n t a l   t e c k e n . 
 ?   m a t c h a r   e x a k t   e t t   t e c k e n . 
 [ a b c ]   m a t c h a r   e t t   t e c k e n   f r � n   u p p s � t t n i n g e n . 
 [ a - z ]   m a t c h a r   e t t   t e c k e n   i   i n t e r v a l l e t . 
 E x e m p e l :   * . h t m l ;   p h o t o ? ? . p n g > M a s k   k a n   u t � k a s   m e d   s � k v � g s m a s k . 
 E x e m p e l :   * / p u b l i c _ h t m l / * . h t m l %M � n s t e r : 
 ! !   u t � k a s   t i l l   u t r o p s t e c k e n 
 !   u t � k a s   t i l l   f i l n a m n 
 ! &   u t � k a s   t i l l   l i s t a   m e d   v a l d a   f i l e r   ( c i t a t ,   s p a c e - a v g r � n s a t ) 
 ! /   u t � k a s   t i l l   a k t u e l l   f j � r r s � k v � g 
 ! @   u t � k a s   t i l l   a k t u e l l   s e s s i o n s v � r d n a m n 
 ! U   u t � k a s   t i l l   a k t u e l l   s e s s i o n s a n v � n d a r n a m n 
 ! P   u t � k a s   t i l l   a k t u e l l   s e s s i o n s l � s e n o r d 
 ! ? p r o m p t [ \ ] ? s t a n d a r d !   u t � k a s   t i l l   a n v � n d a r d e f i n i e r a t   v � r d e   m e d   g i v e n   p r o m p t   o c h   s t a n d a r d   ( a l t e r n a t i v   \   u n d v i k e r   e s c a p e ) 
 ! ` c o m m a n d `   u t � k a s   t i l l   o u t p u t   a v   l o k a l t   k o m m a n d o 
   
 L o k a l t   m � n s t e r k o m m a n d o : 
 ! ^ !   u t � k a s   t i l l   f i l n a m n   f r � n   l o k a l   p a n e l 
   
 E x e m p e l : 
 g r e p   " ! ? M � n s t e r : ? ! "   ! & A A l l a   � v e r f � r i n g a r   i   b a k g r u n d e n   s l u t f � r d e s .   A n s l u t n i n g   a v s l u t a d e s .   L � s n i n g   a v   f j � r r k a t a l o g   a v b r � t s . ( S y n k r o n i s e r a d   b l � d d r i n g   s a t t e s   % s . | p � | a v ' V i s n i n g   a v   d o l d a   f i l e r   s a t t e s   % s . | p � | a v G A u t o m a t i s k   u p p d a t e r i n g   a v   f j � r r k a t a l o g   e f t e r   o p e r a t i o n   s a t t e s   % s . | p � | a v 1 � v e r f � r i n g   i   b a k g r u n d e n   k r � v e r   d i n   u p p m � r k s a m h e t .  � v e r f � r i n g s k � n   � r   t o m . Z ! Y   � r 
 ! M   m � n a d 
 ! D   d a g 
 ! T   t i d 
 ! P   p r o c e s s   i d 
 ! @   v � r d n a m n 
 ! S   s e s s i o n s n a m n 
 E x e m p e l : C : \ ! S ! T . l o g K P a s s i v t   l � g e   m � s t e   v a r a   a k t i v e r a d   n � r   F T P   a n s l u t n i n g   g e n o m   p r o x y   h a r   v a l t s . L U p p d a t e r i n g s k o n t r o l l   f � r   a p p l i k a t i o n e n   � r   t e m p o r � r t   a v s t � n g d .   F � r s � k   s e n a r e .  & G �   t i l l  V a d   � r   n y t t    O p e r a t i o n e n   s l u t f � r d e s  & P r i n t  & A s s o c i e r a d   a p p l i k a t i o n  P �  A v  A u t o V * * H u v u d l � s e n o r d e t   h a r   � n d r a t s . * * 
 
 D i n a   l a g r a d e   l � s e n o r d   � r   s � k r a d e   m e d   A E S - k r y p t e r i n g .  H u v u d l � s e n o r d e t   h a r   � n d r a t s . S * * D u   h a r   t a g i t   b o r t   h u v u d l � s e n o r d e t . * * 
 
 D i n a   l a g r a d e   l � s e n o r d   � r   i n t e   s � k r a   l � n g r e .  H u v u d l � s e n o r d :    S e n a s t   k o n t r o l l e r a d :   % s  K o m m e r   a t t   k o n t r o l l e r a   i g e n :   % s  S e n a s t e   s e s s i o n e r Q M a s k e r   s k i l j s   � t   m e d   s e m i k o l o n   e l l e r   k o m m a .   
 P l a c e r a   u t e s l u t n a   m a s k e r   e f t e r   p i p e . , M a s k s l u t   m e d   s n e d s t r e c k   v � l j e r   u t   k a t a l o g e r .   � > s t o r l e k   m a t c h a r   f i l   s o m   � r   s t � r r e   � n   s t o r l e k 
 < s t o r l e k   m a t c h a r   f i l   m i n d r e   � n   s t o r l e k 
 > y y y y - m m - d d   m a t c h a r   f i l   s o m   � n d r a t s   e f t e r   d e t   d a t u m e t 
 < y y y y - m m - d d   m a t c h a r   f i l   s o m   � n d r a t s   f � r e   d e t   d a t u m e t 
 E x e m p e l :   * . z i p > 1 G ;   < 2 0 1 2 - 0 1 - 2 1  S e   h j � l p   f � r   f l e r   a l t e r n a t i v .  U T F - 8 � * * F � l j a n d e   a n v � n d a r s t a t i s t i k s d a t a   s k i c k a s   a n o n y m t   t i l l   W i n S C P . * * 
 
 U n d e r   t i d e n   k a n   a n n a n   s t a t i s t i k   s a m l a s   i n ,   k o m   g � r n a   t i l l b a k a   s e n a r e   f � r   a t t   k o n t r o l l e r a   e l l e r   k o n s u l t e r a   h j � l p e n . Z D e t   f i n n s   i n g e n   a n v � n d a r s t a t i s t i k   i n s a m l a d   � n n u .   F � r s � k   i g e n   s e n a r e   e l l e r   k o n s u l t e r a   H j � l p  � p p n a   w e b b p l a t s k a t a l o g   ' % s '  � p p n a r   a r b e t s y t a   ' % s '  S e n a s t e   a r b e t s y t o r  M i n   a r b e t s y t a - A r b e t s y t a   ' % s '   k o m m e r   a t t   s p a r a s   a u t o m a t i s k t .  A r b e t s y t a :   % s _ D u   h a r   v a l t   a t t   i n t e   s e   d i a l o g r u t a n   � v e r f � r i n g s a l t e r n a t i v   n � s t a   g � n g .   K l i c k a   h � r   f � r   a t t   � n g r a .  F � r i n s t � l l n i n g a r 	 A v s l u t a d e u % s 
 
 D e t   u p p s t o d   n � g r a   f e l   v i d   k r y p t e r i n g e n   a v   l � s e n o r d   m e d   h j � l p   a v   e t t   n y t t   h u v u d l � s e n o r d   e l l e r   d e k r y p t e r a   l � s e n o r d . � W i n S C P   � r   e n   f r i   S F T P - k l i e n t   o c h   F T P - k l i e n t   f � r   W i n d o w s   m e d   � p p e n   k � l l k o d .   D e s s   h u v u d s a k l i g a   f u n k t i o n   � r   s � k e r   f i l � v e r f � r i n g   m e l l a n   e n   l o k a l   o c h   f j � r r d a t o r .   U t � v e r   d e t t a   e r b j u d e r   W i n S C P   g r u n d l � g g a n d e   f u n k t i o n a l i t e t   f � r   f i l h a n t e r i n g .  W I N _ F O R M S _ S T R I N G S  I n g e n   s e s s i o n s l o g g .  L o g g n i n g   t i l l   f i l   � r   a v s t � n g d . 
 I n g e n   l o g g  S e s s i o n   ' % s '   l o g g  % s   f i l   ' % s '   t i l l   % s :  % s   % d   f i l e r   t i l l   % s :      l o k a l   k a t a l o g  f j � r r k a t a l o g    F l y t t a 	 s l � p p   m � l            T a r   b o r t  S t � l l e r   i n   i n s t � l l n i n g a r  T e m p o r � r   k a t a l o g 
 N y   k a t a l o g     	 A v m a r k e r a  M a r k e r a  % d   f i l  % d   f i l e r 
 % d   k a t a l o g  % d   k a t a l o g e r  % d   s y m b o l i s k   l � n k  % d   s y m b o l i s k a   l � n k a r    % s   E g e n s k a p e r  % s ,   . . .   E g e n s k a p e r  A n g e   g i l t i g t   g r u p p n a m n .  A n g e   g i l t i g t   � g a r n a m n .  T i l l b a k a   t i l l   % s  F r a m � t   t i l l   % s      A n s l u t n i n g s t i d  K o m p r i m e r i n g   ( % s )      I n f o r m a t i o n   o m   v a l d   f i l 7 K o m p r i m e r i n g   ( k l i e n t   ��  s e r v e r :   % s ,   s e r v e r   ��  k l i e n t :   % s )   P � p p n a   s p a r a d   s e s s i o n   ' % s '   ( h � l l   n e r e   S H I F T   f � r   a t t   � p p n a   s e s s i o n   i   n y t t   f � n s t e r )      L i c e n s   f � r   % s                � p p n a   k a t a l o g  H a n t e r a   b o k m � r k e n             
 R a d :   % d / % d 
 K o l u m n :   % d  T e c k e n :   % d   ( 0 x % . 2 x )  � n d r a d  K a n   i n t e   h i t t a   s t r � n g e n   ' % s ' .  T o t a l t   a n t a l   e r s � t t n i n g a r :   % d  G �   t i l l   r a d 
 R a d n u m m e r :  O g i l t i g t   r a d n u m m e r .  R e d i g e r a   l � n k / g e n v � g  L � g g   t i l l   l � n k / g e n v � g  F r � n k o p p l a d .  A n s l u t e r . . .  V � l j   s e s s i o n   ' % s '  L � g g   t i l l   p l a t s p r o f i l  P l a t s p r o f i l n a m n :    F l y t t a   p l a t s p r o f i l  N y t t   k a t a l o g n a m n :  S p a r a   s e s s i o n   s o m  & S p a r a   s e s s i o n   s o m : $ S p a r a   & l � s e n o r d   ( r e k o m m e n d e r a s   i n t e )    K � r   e g e t   k o m m a n d o  K � r   e g e t   k o m m a n d o   ' % s '          K  R 5 % s ,   % d   p t 
 T h e   Q u i c k   B r o w n   F o x   J u m p s   O v e r   T h e   L a z y   D o g  O k � n d  B e r � k n a   k a t a l o g s t o r l e k        A l l m � n n a   i n s t � l l n i n g a r  L a g r a d e   s e s s i o n e r  C a c h a d e   v � r d n y c k l a r  K o n f i g u r a t i o n e n s   I N I - f i l  S l u m p t a l s f r �   f i l  V � l j   l o k a l   k a t a l o g .  F l y t t a r      F l y t t a  H � l l   f j � r r k a t a l o g e n   u p p d a t e r a d % B e h � l l e r   f j � r r k a t a l o g e n   u p p d a t e r a d . . .    T e m p o r � r a   k a t a l o g e r  N y   f i l  R e d i g e r a   f i l  & S k r i v   f i l n a m n : ( D u p l i c a t e   f i l e   ' % s '   t o   r e m o t e   d i r e c t o r y : ' D u p l i c a t e   % d   f i l e s   t o   r e m o t e   d i r e c t o r y :  D u b b l e r a  K o p i e r a r  L � g g   t i l l   e g e t   k o m m a n d o  R e d i g e r a   e g e t   k o m m a n d o  L  F          H � & m t a   f l e r . . .  V � l j   e d i t o r a p p l i k a t i o n . 0 K � r b a r a   f i l e r   ( * . e x e ) | * . e x e | A l l a   f i l e r   ( * . * ) | * . *  % s   a v   % s   i   % s   a v   % s , L � g g   t i l l   f � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g + R e d i g e r a   f � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g 	 S & t a n d a r d  & K o n f i g u r e r a . . .  E g & e t . . .  E g e t   k o m m a n d o  L � g g   t i l l   e d i t o r  R e d i g e r a   e d i t o r  % s ,   B a s e r a s   p �   % s   v e r s i o n   % s  & � p p n a  & K o p i e r a  E n d a s t   & s a m m a   s t o r l e k   N u m b e r   o f   L i c e n s e s :   % s | U n l i m i t e d  P r o d u c t   I D :   % s  % s   ( E x p i r a t i o n   o n   % s )  % s       E d u c a t i o n a l   L i c e n s e  H � m t a r   e g e n s k a p e r    S S H   i m p l e m e n t a t i o n  K r y p t e r i n g s a l g o r i t m  K o m p r i m e r i n g  F i l � v e r f � r i n g s p r o t o k o l l  K a n   � n d r a   r � t t i g h e t e r  K a n   � n d r a   � g a r e / g r u p p  K a n   k � r a   g o d t y c k l i g t   k o m m a n d o " K a n   s k a p a   s y m b o l i s k   l � n k / h � r d   l � n k  K a n   s l �   u p p   a n v � n d a r g r u p p e r  K a n   d u b b l e r a   f j � r r f i l e r   $ � v e r f � r i n g s l � g e   f � r   r e n   t e x t   ( A S C I I ) $ K a n   k o n t r o l l e r a   t i l l g � n g l i g t   u t r y m m e  T o t a l t   a n t a l   b y t e s   p �   e n h e t  L e d i g t   a n t a l   b y t e s   p �   e n h e t   T o t a l t   a n t a l   b y t e s   f � r   a n v � n d a r e  L e d i g a   b y t e s   f � r   a n v � n d a r e  B y t e s   p e r   a l l o k e r i n g s e n h e t  O k � n d " H i t t a   P u T T Y / T e r m i n a l k l i e n t   k � r b a r a P P u T T Y / T e r m i n a l k l i e n t   k � r b a r a | % s | K � r b a r a   f i l e r   ( * . e x e ) | * . e x e | A l l a   f i l e r   ( * . * ) | * . *  % s   a v   % s | N / A  J � m f � r  S y n k r o n i s e r i n g  A u t e n t i s e r i n g s b a n e r * I N I - f i l   ( * . i n i ) | * . i n i | A l l a   f i l e r   ( * . * ) | * . * ) V � l j   f i l   a t t   e x p o r t e r a   i n s t � l l n i n g a r   t i l l    S & e n a s t e :   % s  S & e n a s t e  B e r � k n a r   f i l k o n t r o l l s u m m a  K a n   b e r � k n a   f i l k o n t r o l l s u m m a  O k � n d  P r o t o k o l l   s o m   a n v � n d s    O s � k e r   a n s l u t n i n g  S � k e r   a n s l u t n i n g   ( % s )  E n d a s t   p r o t o k o l l k o m m a n d o n  F j � r r s y s t e m  K r y p t o g r a f i s k t   p r o t o k o l l      M i n a   d o k u m e n t 	 S k r i v b o r d    K o m m a n d o  S � t t   t i l l   s & t a n d a r d  - -   v a r n a   e f t e r   d e t t a   - -  3 D E S  B l o w f i s h  A E S   ( e n d a s t   S S H - 2 )  D E S  A r c f o u r   ( e n d a s t   S S H - 2 )  - -   v a r n a   e f t e r   d e t t a   - -  D i f f i e - H e l l m a n   g r u p p   1  D i f f i e - H e l l m a n   g r u p p   1 4  D i f f i e - H e l l m a n   g r u p p   u t b y t e  R S A - b a s e r a t   n y c k e l u t b y t e      V � l j   l o k a l   p r o x y a p p l i k a t i o n   � M � n s t e r : 
 \ n   f � r   n y   r a d 
 \ r   f � r   v a g n r e t u r 
 \ t   f � r   t a b 
 \ x X X   f � r   h e x a d e c i m a l   a s c i i k o d 
 \ \   f � r   b a c k s l a s h 
 % v � r d   u t � k a s   t i l l   v � r d n a m n 
 % p o r t   u t � k a s   t i l l   p o r t n u m m e r 
 % u a n v � n d a r e   u t � k a s   t i l l   p r o x y a n v � n d a r n a m n 
 % l � s e n   u t � k a s   t i l l   p r o x y l � s e n o r d 
 % %   f � r   p r o c e n t t e c k e n = W e b b p l a t s k a t a l o g   e l l e r   a r b e t s y t a   m e d   n a m n e t   ' % s '   f i n n s   r e d a n . E � r   d u   s � k e r   a t t   d u   v i l l   r a d e r a   s e s s i o n s k a t a l o g   ' % s '   m e d   % d   s e s s i o n e r ? $ K a n   i n t e   r a d e r a   s p e c i a l s e s s i o n   ' % s ' .  S k a p a   s e s s i o n s k a t a l o g  N y t t   k a t a l o g n a m n : ! � p p n a   s p a r a d   s e s s i o n s k a t a l o g   ' % s '  H o w   t o   p u r c h a s e   a   l i c e n s e . . .  M � l & k a t a l o g : � * * V i l l   d u   � p p n a   e n   s e p a r a t   s k a l s e s s i o n   f � r   a t t   d u b b l e r a   f i l e n ? * * 
 
 A k t u e l l   s e s s i o n   s t � d e r   i n t e   d i r e k t   d u b b l e r i n g   a v   f j � r r f i l e r .   S e p a r a t a   s k a l s e s s i o n e r   k a n   � p p n a s   f � r   a t t   b e a r b e t a   d u b b l e r i n g e n .   A l t e r n a t i v t   k a n   d u   d u b b l e r a   f i l e n   v i a   e n   l o k a l   t e m p o r � r   k o p i a .  E d i t o r  % s   ( % s )  % d   d o l d  % d   f i l t r e r a s  F i l t e r � A k t u e l l   s e s s i o n   t i l l � t e r   e n d a s t   f � r � n d r i n g   a v   U I D   � g a n d e t .   D e t   v a r   i n t e   m � j l i g t   a t t   l � s a   U I D   f r � n   k o n t o n a m n e t   " % s " .   S p e c i f i c e r a   U I D   e x p l i c i t   i s t � l l e t .  � v e r f � r   i   & b a k g r u n d e n  % s   ( l � g g   t i l l   i   � v e r f � r i n g s k � )  I n g e n  V � l j   k o r t k o m m a n d o  K o r & t k o m m a n d o : 
 O b e g r � n s a t  H u v u d l � s e n o r d  & N u v a r a n d e   h u v u d l � s e n o r d :  N & y t t   h u v u d l � s e n o r d :  U p p r e p a   h u v u d l � s e n o r d : - S p a r a   & l � s e n o r d   ( s k y d d a s   g e n o m   h u v u d l � s e n o r d ) 	 L e t a   i   % s  S � k 	 S � k e r   . . .  K l a r . 	 A v b r u t e n .    & S t a r t  & S t o p p  S p a r a   & l � s e n o r d  A v b r y t e r . . .  K o d n i n g :   % s c F i l e n   h a r   � n d r a t s .   � n d r i n g a r   k o m m e r   a t t   g �   f � r l o r a d e ,   o m   f i l e n   l a d d a s   m e d   a n n a n   k o d n i n g .   F o r t s � t t a ? F � r   d u   s � k e r   p �   a t t   d u   v i l l   t a   b o r t   a r b e t s y t a n   ' % s '   m e d   % d   s e s s i o n ( e r ) ?    S p a r a   a r b e t s y t a   s o m  & S p a r a   a r b e t s y t a   s o m : $ S p a r a   & l � s e n o r d   ( r e k o m m e n d e r a s   i n t e ) . S p a r a   & l � s e n o r d   ( s o m   s k y d d a s   a v   h u v u d l � s e n o r d )  S p a r a   & l � s e n o r d Q � p p n a   a r b e t s y t a   ' % s '   ( h � l l   n e r   S h i f t   f � r   a t t   � p p n a   a r b e t s y t a n   i   e t t   n y t t   f � n s t e r )  & � p p n a   k a t a l o g U � p p n a   w e b b p l a t s k a t a l o g   ' % s '   ( h � l l   n e r   S h i f t   f � r   a t t   � p p n a   k a t a l o g   i   e t t   n y t t   f � n s t e r )    & S k a p a   g e n v � g   p �   s k r i v b o r d e t , A k t i v e r a   & a u t o m a t i s k t   s p a r a n d e   a v   a r b e t s y t a n  H � m t a  � v e r f � r  H � m t a  � v e r f � r ) % s   f i l   ' % s '   t i l l   % s   o c h   t a   b o r t   o r i g i n a l : + % s   % d   f i l e r   t i l l   % s   o c h   t a   b o r t   o r i g i n a l e n :  H � m t a   o c h   t a   b o r t  � v e r f � r   o c h   t a   b o r t  K �  I m p o r t e r a   w e b b p l a t s e r - F e l   v i d   l a d d n i n g   a v   f i l   ' % s '   m e d   ' % s '   k o d n i n g                        F e l   v i d   l a d d n i n g   a v   f i l   ' % s ' .  � t e r g � r   t i l l   ' % s '   k o d n i n g . ) V � l j   f i l   a t t   i m p o r t e r a   k o n f i g u r a t i o n   f r � n  S � k :   % s  ( t r y c k   p �   T a b   f � r   n � s t a )  � v e r f � r  H � m t a r  % d   i   k �   �M � n s t e r : 
 ! !   e x p a n d e r a r   t i l l   u t r o p s t e c k e n 
 ! /   e x p a n d e r a r   t i l l   a k t u e l l   f j � r r s � k v � g 
 ! @   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s   v � r d n a m n 
 ! U   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s   a n v � n d a r n a m n 
 ! P   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s   l � s e n o r d 
 ! ? p r o m p t [ \ ] ? d e f a u l t !   e x p a n d e r a r   t i l l   a n v � n d a r v a l t   v � r d e   m e d   g i v e n   p r o m p t   o c h   s t a n d a r d   ( a l t e r n a t i v t   \   u n d v i k e r   e s c a p e ) 
 ! ` c o m m a n d `   e x p a n d e r a r   t i l l   u t d a t a   a v   l o k a l t   k o m m a n d o  N y   w e b b p l a t s  K a t a l o g   w e b b p l a t s 	 A r b e t s y t a D D e t t a   k o m m e r   a t t   a v b r y t a   r e d i g e r i n g   a v   w e b b p l a t s .   V i l l   d u   f o r t s � t t a ? 	 & K a t a l o g :  < r o o t >  S k a l  S C P / S k a l  E d i t o r  & I n g e n   f � r g 2 � t e r s t � l l   s e s s i o n   ( p a n e l )   f � r g   t i l l   s y s t e m s t a n d a r d  F & l e r   f � r g e r . . .  V � l j   f � r g   p �   s e s s i o n   ( p a n e l )      A n s l u t e n 0 A n s l u t e n   m e d   % s .   V � n t a r   p �   v � l k o m s t m e d d e l a n d e . . .   * A n s l u t e n   m e d   % s ,   f � r m e d l a r   S S L - k o p p l i n g . . .  A n s l u t e r   t i l l   % s   . . .  L i s t n i n g   a v   k a t a l o g e r   l y c k a d  K o p p l a r   i f r � n   s e r v e r    s t a r t a r   n e r l a d d n i n g   a v   % s  N e r l a d d n i n g   l y c k a d   * F � r s � k e r   a t t   a n s l u t a   % s   g e n o m   F T P   p r o x y . . .                 � t e r f � r   l i s t n i n g   a v   k a t a l o g e r . . . 7 S S L - k o p p l i n g   u p p r � t t a d .   V � n t a r   p �   v � l k o m s t m e d d e l a n d e . . .  S S L - k o p p l i n g   u p p r � t t a d  S t a r t a r   � v e r f � r i n g   a v   % s  � v e r f � r i n g   l y c k a d     # H � m t a r   f i l i n f o r m a t i o n   f r a m g � n g s r i k t  H � m t a r   f i l i n f o r m a t i o n . . .  K u n d e   i n t e   h � m t a   f i l i n f o r m a t i o n                   5 K u n d e   i n t e   s k a p a   s o c k e t   i   d e n   a n g i v n a   p o r t i n t e r v a l l e t    K a n   i n t e   u p p r � t t a   S S L - k o p p l i n g   ' K u n d e   i n t e   � t e r f �   l i s t n i n g   a v   k a t a l o g e r     # K a n   i n t e   i n i t i a l i s e r a   S S L - b i b l i o t e k         , � v e r f � r i n g s t u n n e l   k a n   i n t e   � p p n a s .   O r s a k :   % s    K a n   i n t e   t o l k a   v � r d n a m n   " % s " > � t e r u p p t a g n i n g s k o m m a n d o   s t � d s   i n t e   a v   s e r v e r ,   s k r i v a   � v e r   f i l . I P a u s k o m m a n d o   s t � d s   i n t e   a v   s e r v e r ,   m e n   l o k a l   o c h   f j � r r f i l s t o r l e k   � r   l i k a . , O f � r m � g e n   a t t   s k i c k a   k o m m a n d o .   K o p p l a   i f r � n .    P e e r   c e r t i f i k a t   f � r k a s t a s    N e r l a d d n i n g   a v b r u t e n                      F i l e n   f i n n s   r e d a n          P r o x y   k r � v e r   a u t e n t i s e r i n g P N � d v � n d i g   a u t e n t i s e r i n g s t y p   r a p p o r t e r a d   a v   p r o x y s e r v e r   � r   o k � n d   e l l e r   s t � d s   i n t e % K a n   i n t e   a v g � r a   v � r d   t i l l   p r o x y s e r v e r ! K a n   i n t e   a n s l u t a   t i l l   p r o x y s e r v e r C B e g � r a n   f r � n   p r o x y   m i s s l y c k a d e s ,   k a n   i n t e   a n s l u t a   g e n o m   p r o x y s e r v e r                        T i m e o u t   d e t e k t e r a d .  � v e r f � r i n g   a v b r u t e n            K u n d e   i n t e   s � t t a   f i l p e k a r e  O k � n t   f e l   i   S S L - l a g r e t % K u n d e   i n t e   v e r i f i e r a   S S L - c e r t i f i k a t e t                                               1 � v e r s � t t n i n g :   A .   P e t t e r s s o n   < a z @ k t h . s e >   2 0 0 8 - 2 0 1 4                W I N _ V A R I A B L E $ C o p y r i g h t   �   2 0 0 0 - 2 0 1 4   M a r t i n   P r i k r y l  h t t p : / / w i n s c p . n e t / " h t t p : / / w i n s c p . n e t / e n g / d o c s / h i s t o r y    h t t p : / / w i n s c p . n e t / f o r u m /  h t t p : / / w i n s c p . n e t / u p d a t e s . p h p " h t t p : / / w i n s c p . n e t / e n g / d o w n l o a d . p h p   h t t p : / / w i n s c p . n e t / e n g / d o n a t e . p h p * h t t p : / / w i n s c p . n e t / e n g / d o c s / ? v e r = % s & l a n g = % s , h t t p : / / w i n s c p . n e t / e n g / d o c s / % s ? v e r = % s & l a n g = % s & h t t p : / / w i n s c p . n e t / e n g / t r a n s l a t i o n s . p h p 9 h t t p : / / w i n s c p . n e t / e n g / d o c s / s e a r c h . p h p ? q = % s & v e r = % s & l a n g = % s N h t t p : / / w i n s c p . n e t / f o r u m / p o s t i n g . p h p ? m o d e = n e w t o p i c & f = 2 & r e p o r t = % s & v e r = % s & l a n g = % s ! h t t p : / / w i n s c p . n e t / e n g / u p g r a d e . p h p                  a n   u n n a m e d   f i l e                      N o   e r r o r   m e s s a g e   i s   a v a i l a b l e . ' A n   u n s u p p o r t e d   o p e r a t i o n   w a s   a t t e m p t e d . $ A   r e q u i r e d   r e s o u r c e   w a s   u n a v a i l a b l e .  O u t   o f   m e m o r y .  A n   u n k n o w n   e r r o r   h a s   o c c u r r e d .                                        F a i l e d   t o   l a u n c h   h e l p .  I n t e r n a l   a p p l i c a t i o n   e r r o r .  C o m m a n d   f a i l e d . ) I n s u f f i c i e n t   m e m o r y   t o   p e r f o r m   o p e r a t i o n . P S y s t e m   r e g i s t r y   e n t r i e s   h a v e   b e e n   r e m o v e d   a n d   t h e   I N I   f i l e   ( i f   a n y )   w a s   d e l e t e d . B N o t   a l l   o f   t h e   s y s t e m   r e g i s t r y   e n t r i e s   ( o r   I N I   f i l e )   w e r e   r e m o v e d . F T h i s   p r o g r a m   r e q u i r e s   t h e   f i l e   % s ,   w h i c h   w a s   n o t   f o u n d   o n   t h i s   s y s t e m . t T h i s   p r o g r a m   i s   l i n k e d   t o   t h e   m i s s i n g   e x p o r t   % s   i n   t h e   f i l e   % s .   T h i s   m a c h i n e   m a y   h a v e   a n   i n c o m p a t i b l e   v e r s i o n   o f   % s .      P l e a s e   e n t e r   a n   i n t e g e r .  P l e a s e   e n t e r   a   n u m b e r . * P l e a s e   e n t e r   a n   i n t e g e r   b e t w e e n   % 1   a n d   % 2 . ( P l e a s e   e n t e r   a   n u m b e r   b e t w e e n   % 1   a n d   % 2 . ( P l e a s e   e n t e r   n o   m o r e   t h a n   % 1   c h a r a c t e r s .  P l e a s e   s e l e c t   a   b u t t o n . * P l e a s e   e n t e r   a n   i n t e g e r   b e t w e e n   0   a n d   2 5 5 .   P l e a s e   e n t e r   a   p o s i t i v e   i n t e g e r .   P l e a s e   e n t e r   a   d a t e   a n d / o r   t i m e .  P l e a s e   e n t e r   a   c u r r e n c y .                U n e x p e c t e d   f i l e   f o r m a t . V % 1 
 C a n n o t   f i n d   t h i s   f i l e . 
 P l e a s e   v e r i f y   t h a t   t h e   c o r r e c t   p a t h   a n d   f i l e   n a m e   a r e   g i v e n .  D e s t i n a t i o n   d i s k   d r i v e   i s   f u l l . 5 U n a b l e   t o   r e a d   f r o m   % 1 ,   i t   i s   o p e n e d   b y   s o m e o n e   e l s e . A U n a b l e   t o   w r i t e   t o   % 1 ,   i t   i s   r e a d - o n l y   o r   o p e n e d   b y   s o m e o n e   e l s e . . A n   u n e x p e c t e d   e r r o r   o c c u r r e d   w h i l e   r e a d i n g   % 1 . . A n   u n e x p e c t e d   e r r o r   o c c u r r e d   w h i l e   w r i t i n g   % 1 .                                           # U n a b l e   t o   r e a d   w r i t e - o n l y   p r o p e r t y . # U n a b l e   t o   w r i t e   r e a d - o n l y   p r o p e r t y .      N o   e r r o r   o c c u r r e d . - A n   u n k n o w n   e r r o r   o c c u r r e d   w h i l e   a c c e s s i n g   % 1 .  % 1   w a s   n o t   f o u n d .  % 1   c o n t a i n s   a n   i n v a l i d   p a t h . = % 1   c o u l d   n o t   b e   o p e n e d   b e c a u s e   t h e r e   a r e   t o o   m a n y   o p e n   f i l e s .  A c c e s s   t o   % 1   w a s   d e n i e d . . A n   i n v a l i d   f i l e   h a n d l e   w a s   a s s o c i a t e d   w i t h   % 1 . < % 1   c o u l d   n o t   b e   r e m o v e d   b e c a u s e   i t   i s   t h e   c u r r e n t   d i r e c t o r y . 6 % 1   c o u l d   n o t   b e   c r e a t e d   b e c a u s e   t h e   d i r e c t o r y   i s   f u l l .  S e e k   f a i l e d   o n   % 1 5 A   h a r d w a r e   I / O   e r r o r   w a s   r e p o r t e d   w h i l e   a c c e s s i n g   % 1 . 0 A   s h a r i n g   v i o l a t i o n   o c c u r r e d   w h i l e   a c c e s s i n g   % 1 . 0 A   l o c k i n g   v i o l a t i o n   o c c u r r e d   w h i l e   a c c e s s i n g   % 1 .  D i s k   f u l l   w h i l e   a c c e s s i n g   % 1 . . A n   a t t e m p t   w a s   m a d e   t o   a c c e s s   % 1   p a s t   i t s   e n d .    N o   e r r o r   o c c u r r e d . - A n   u n k n o w n   e r r o r   o c c u r r e d   w h i l e   a c c e s s i n g   % 1 . / A n   a t t e m p t   w a s   m a d e   t o   w r i t e   t o   t h e   r e a d i n g   % 1 . . A n   a t t e m p t   w a s   m a d e   t o   a c c e s s   % 1   p a s t   i t s   e n d . 0 A n   a t t e m p t   w a s   m a d e   t o   r e a d   f r o m   t h e   w r i t i n g   % 1 .  % 1   h a s   a   b a d   f o r m a t . " % 1   c o n t a i n e d   a n   u n e x p e c t e d   o b j e c t .   % 1   c o n t a i n s   a n   i n c o r r e c t   s c h e m a .                 � S e t t i n g   b i t   t r a n s p a r e n c y   c o l o r   i s   n o t   a l l o w e d   f o r   p n g   i m a g e s   c o n t a i n i n g   a l p h a   v a l u e   f o r   e a c h   p i x e l   ( C O L O R _ R G B A L P H A   a n d   C O L O R _ G R A Y S C A L E A L P H A ) O T h i s   o p e r a t i o n   i s   n o t   v a l i d   b e c a u s e   t h e   c u r r e n t   i m a g e   c o n t a i n s   n o   v a l i d   h e a d e r . 4 T h e   n e w   s i z e   p r o v i d e d   f o r   i m a g e   r e s i z i n g   i s   i n v a l i d . o T h e   " P o r t a b l e   N e t w o r k   G r a p h i c s "   c o u l d   n o t   b e   c r e a t e d   b e c a u s e   i n v a l i d   i m a g e   t y p e   p a r a m e t e r s   h a v e   b e i n g   p r o v i d e d .                         [ C o u l d   n o t   d e c o m p r e s s   t h e   i m a g e   b e c a u s e   i t   c o n t a i n s   i n v a l i d   c o m p r e s s e d   d a t a .  
   D e s c r i p t i o n :   B T h e   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   c o n t a i n s   a n   i n v a l i d   p a l e t t e . � T h e   f i l e   b e i n g   r e a d   i s   n o t   a   v a l i d   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   b e c a u s e   i t   c o n t a i n s   a n   i n v a l i d   h e a d e r .   T h i s   f i l e   m a y   b e   c o r r u p t e d ,   t r y   o b t a i n i n g   i t   a g a i n n T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   n o t   s u p p o r t e d   o r   i t   m i g h t   b e   i n v a l i d .  
 ( I H D R   c h u n k   i s   n o t   t h e   f i r s t ) � T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   n o t   s u p p o r t e d   b e c a u s e   e i t h e r   i t s   w i d t h   o r   h e i g h t   e x c e e d s   t h e   m a x i m u m   s i z e   o f   6 5 5 3 5   p i x e l s .  T h e r e   i s   n o   s u c h   p a l e t t e   e n t r y . d T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   c o n t a i n s   a n   u n k n o w n   c r i t i c a l   p a r t   w h i c h   c o u l d   n o t   b e   d e c o d e d . p T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   e n c o d e d   w i t h   a n   u n k n o w n   c o m p r e s s i o n   s c h e m e   w h i c h   c o u l d   n o t   b e   d e c o d e d . c T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   u s e s   a n   u n k n o w n   i n t e r l a c e   s c h e m e   w h i c h   c o u l d   n o t   b e   d e c o d e d . - T h e   c h u n k s   m u s t   b e   c o m p a t i b l e   t o   b e   a s s i g n e d . j T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   i n v a l i d   b e c a u s e   t h e   d e c o d e r   f o u n d   a n   u n e x p e c t e d   e n d   o f   t h e   f i l e . 8 T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   c o n t a i n s   n o   d a t a . ] T h e   p r o g r a m   t r i e d   t o   a d d   a   e x i s t e n t   c r i t i c a l   c h u n k   t o   t h e   c u r r e n t   i m a g e   w h i c h   i s   n o t   a l l o w e d . I I t ' s   n o t   a l l o w e d   t o   a d d   a   n e w   c h u n k   b e c a u s e   t h e   c u r r e n t   i m a g e   i s   i n v a l i d . 7 T h e   p n g   i m a g e   c o u l d   n o t   b e   l o a d e d   f r o m   t h e   r e s o u r c e   I D . o S o m e   o p e r a t i o n   c o u l d   n o t   b e   p e r f o r m e d   b e c a u s e   t h e   s y s t e m   i s   o u t   o f   r e s o u r c e s .   C l o s e   s o m e   w i n d o w s   a n d   t r y   a g a i n .  N o   a c t i v e   d o c u m e n t  N o d e   " % s "   n o t   f o u n d  I D O M N o d e   r e q u i r e d . A t t r i b u t e s   a r e   n o t   s u p p o r t e d   o n   t h i s   n o d e   t y p e  I n v a l i d   n o d e   t y p e + M i s m a t c h e d   p a r a m a t e r s   t o   R e g i s t e r C h i l d N o d e s 0 E l e m e n t   " % s "   d o e s   n o t   c o n t a i n   a   s i n g l e   t e x t   n o d e 4 D O M   I m p l e m e n t a t i o n   d o e s   n o t   s u p p o r t   I D O M P a r s e O p t i o n s # I t e m T a g   p r o p e r t y   i s   n o t   i n i t i a l i z e d  N o d e   i s   r e a d o n l y C R e f r e s h   i s   o n l y   s u p p o r t e d   i f   t h e   F i l e N a m e   o r   X M L   p r o p e r t i e s   a r e   s e t  F i l e N a m e   c a n n o t   b e   b l a n k  L i n e j T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   n o t   v a l i d   b e c a u s e   i t   c o n t a i n s   i n v a l i d   p i e c e s   o f   d a t a   ( c r c   e r r o r ) y T h e   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   c o u l d   n o t   b e   l o a d e d   b e c a u s e   o n e   o f   i t s   m a i n   p i e c e   o f   d a t a   ( i h d r )   m i g h t   b e   c o r r u p t e d U T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   i n v a l i d   b e c a u s e   i t   h a s   m i s s i n g   i m a g e   p a r t s .  & S k a p a   g e n v � g   h i t  & A v b r y t  T o o l b a r   i t e m   i n d e x   o u t   o f   r a n g e  T o o l b a r   i t e m   a l r e a d y   i n s e r t e d ? A n   i t e m   v i e w e r   a s s o c i a t e d   t h e   s p e c i f i e d   i t e m   c o u l d   n o t   b e   f o u n d  M o r e   B u t t o n s | J A   T T B D o c k   c o n t r o l   c a n n o t   b e   p l a c e d   i n s i d e   a   t o o l   w i n d o w   o r   a n o t h e r   T T B D o c k C C a n n o t   c h a n g e   P o s i t i o n   o f   a   T T B D o c k   i f   i t   a l r e a d y   c o n t a i n s   c o n t r o l s G C a n n o t   s a v e   d o c k a b l e   w i n d o w ' s   p o s i t i o n   b e c a u s e   N a m e   p r o p e r t y   i s   n o t   s e t O C a n n o t   s a v e   d o c k a b l e   w i n d o w ' s   p o s i t i o n   b e c a u s e   D o c k e d T o ' s   N a m e   p r o p e r t y   n o t   s e t ) " % s "   D O M I m p l e m e n t a t i o n   a l r e a d y   r e g i s t e r e d  N o   m a t c h i n g   D O M   V e n d o r :   " % s " < S e l e c t e d   D O M   V e n d o r   d o e s   n o t   s u p p o r t   t h i s   p r o p e r t y   o r   m e t h o d ; P r o p e r t y   o r   M e t h o d   " % s "   i s   n o t   s u p p o r t e d   b y   D O M   V e n d o r   " % s "  N o d e   c a n n o t   b e   n u l l   M i c r o s o f t   M S X M L   i s   n o t   i n s t a l l e d  � n d r a d  A t t r  E x t  F i l e s y s t e m   O p e r a t i o n 	 \ / : * ? " < > |    ' N e w   n a m e   c o n t a i n s   i n v a l i d   c h a r a c t e r s   % s  F i l o p e r a t i o n  % s   � r   e n   o g i l t i g   e n h e t s b o k s t a v .  R � t t i g h e t e r  � g a r e  G r u p p  M � l   l � n k  F i l t y p  & K o p i e r a   h i t  & F l y t t a   h i t    F i l e n   f i n n s   r e d a n :   % F i l n a m n e t   i n n e h � l l e r   o g i l t i g a   t e c k e n :  F i l   % s  % u   F i l e r  % u   K a t a l o g e r  H u v u d k a t a l o g * K a n   i n t e   a v s l u t a   t r � d   f � r   i k o n u p p d a t e r i n g .  D r a S l � p p   f e l :   % d  E n h e t   ' % s : '   � r   i n t e   k l a r .  K a t a l o g e n   ' % s '   f i n n s   i n t e .  D r a g & d r o p   e r r o r :   % d  /   < r o o t >  F i l s y s t e m s o p e r a t i o n  N a m n  S t o r l e k  F i l t y p  S t a r t   i n d e x   o u t   o f   b o u n d s   ( % d )  I n v a l i d   c o u n t   ( % d )  I n v a l i d   d e s t i n a t i o n   i n d e x   ( % d )  I n v a l i d   c o d e   p a g e  I n v a l i d   e n c o d i n g   n a m e  B l � d d r a  A l l a   f i l e r   ( * . * ) | * . *  O g i l t i g t   f i l n a m n   -   % s  S o c k e t   e r r o r   ( % s )  T i m e o u t 	 O k � n t   f e l  R e c e i v e d   r e s p o n s e   % d   % s   f r o m   % s " E x c e e d e d   m a x i m a l   r e d i r e c t   l i m i e   % d # K a n   i n t e   h i t t a   n � g o n   g i l t i g   s � k v � g .  U N C   s � k v � g a r   s t � d s   i n t e . ) K a n   i n t e   b y t a   n a m n   p �   f i l   e l l e r   k a t a l o g :    T u e  W e d  T h u  F r i  S a t  S u n d a y  M o n d a y  T u e s d a y 	 W e d n e s d a y  T h u r s d a y  F r i d a y  S a t u r d a y  U n a b l e   t o   c r e a t e   d i r e c t o r y  I n v a l i d   s o u r c e   a r r a y  I n v a l i d   d e s t i n a t i o n   a r r a y " C h a r a c t e r   i n d e x   o u t   o f   b o u n d s   ( % d )  N o v  D e c  J a n u a r y  F e b r u a r y  M a r c h  A p r i l  M a y  J u n e  J u l y  A u g u s t 	 S e p t e m b e r  O c t o b e r  N o v e m b e r  D e c e m b e r  S u n  M o n  F e a t u r e   n o t   i m p l e m e n t e d  % s   ( % s ,   l i n e   % d )  A b s t r a c t   E r r o r ? A c c e s s   v i o l a t i o n   a t   a d d r e s s   % p   i n   m o d u l e   ' % s ' .   % s   o f   a d d r e s s   % p  S y s t e m f e l .     K o d :   % d .  
 % s * E t t   a n r o p   t i l l   e n   O S   f u n k t i o n   m i s s l y c k a d e s  J a n  F e b  M a r  A p r  M a y  J u n  J u l  A u g  S e p  O c t / C u s t o m   v a r i a n t   t y p e   ( % s % . 4 x )   a l r e a d y   u s e d   b y   % s * C u s t o m   v a r i a n t   t y p e   ( % s % . 4 x )   i s   n o t   u s a b l e 2 T o o   m a n y   c u s t o m   v a r i a n t   t y p e s   h a v e   b e e n   r e g i s t e r e d 5 C o u l d   n o t   c o n v e r t   v a r i a n t   o f   t y p e   ( % s )   i n t o   t y p e   ( % s ) = O v e r f l o w   w h i l e   c o n v e r t i n g   v a r i a n t   o f   t y p e   ( % s )   i n t o   t y p e   ( % s )  V a r i a n t   o v e r f l o w  I n v a l i d   a r g u m e n t  I n v a l i d   v a r i a n t   t y p e  O p e r a t i o n   n o t   s u p p o r t e d  U n e x p e c t e d   v a r i a n t   e r r o r  E x t e r n a l   e x c e p t i o n   % x  A s s e r t i o n   f a i l e d  I n t e r f a c e   n o t   s u p p o r t e d  E x c e p t i o n   i n   s a f e c a l l   m e t h o d  O b j e c t   l o c k   n o t   o w n e d ( M o n i t o r   s u p p o r t   f u n c t i o n   n o t   i n i t i a l i z e d   ( E x c e p t i o n   % s   i n   m o d u l e   % s   a t   % p .  
 % s % s  
  A p p l i c a t i o n   E r r o r 1 F o r m a t   ' % s '   i n v a l i d   o r   i n c o m p a t i b l e   w i t h   a r g u m e n t  N o   a r g u m e n t   f o r   f o r m a t   ' % s ' " V a r i a n t   m e t h o d   c a l l s   n o t   s u p p o r t e d  R e a d  W r i t e  F o r m a t   s t r i n g   t o o   l o n g $ E r r o r   c r e a t i n g   v a r i a n t   o r   s a f e   a r r a y ) V a r i a n t   o r   s a f e   a r r a y   i n d e x   o u t   o f   b o u n d s  V a r i a n t   o r   s a f e   a r r a y   i s   l o c k e d  I n v a l i d   v a r i a n t   t y p e   c o n v e r s i o n  I n v a l i d   v a r i a n t   o p e r a t i o n  I n v a l i d   N U L L   v a r i a n t   o p e r a t i o n % I n v a l i d   v a r i a n t   o p e r a t i o n   ( % s % . 8 x ) 
 % s , C u s t o m   v a r i a n t   t y p e   ( % s % . 4 x )   i s   o u t   o f   r a n g e    I n v a l i d   n u m e r i c   i n p u t  D i v i s i o n   b y   z e r o  R a n g e   c h e c k   e r r o r  I n t e g e r   o v e r f l o w   I n v a l i d   f l o a t i n g   p o i n t   o p e r a t i o n  F l o a t i n g   p o i n t   d i v i s i o n   b y   z e r o  F l o a t i n g   p o i n t   o v e r f l o w  F l o a t i n g   p o i n t   u n d e r f l o w  I n v a l i d   p o i n t e r   o p e r a t i o n  I n v a l i d   c l a s s   t y p e c a s t 0 A c c e s s   v i o l a t i o n   a t   a d d r e s s   % p .   % s   o f   a d d r e s s   % p  A c c e s s   v i o l a t i o n  S t a c k   o v e r f l o w  C o n t r o l - C   h i t  P r i v i l e g e d   i n s t r u c t i o n  O p e r a t i o n   a b o r t e d   L C a n n o t   h a v e   m u l t i p l e   s i n g l e   c a s t   o b s e r v e r s   a d d e d   t o   t h e   o b s e r v e r s   c o l l e c t i o n 4 T h e   o b j e c t   d o e s   n o t   i m p l e m e n t   t h e   o b s e r v e r   i n t e r f a c e G N o   s i n g l e   c a s t   o b s e r v e r   w i t h   I D   % s   w a s   a d d e d   t o   t h e   o b s e r v e r   c o l l e c t i o n F N o   m u l t i   c a s t   o b s e r v e r   w i t h   I D   % s   w a s   a d d e d   t o   t h e   o b s e r v e r   c o l l e c t i o n  O b s e r v e r   i s   n o t   a v a i l a b l e 	 < u n k n o w n > ( ' % s '   i s   n o t   a   v a l i d   f l o a t i n g   p o i n t   v a l u e   ' % d . % d '   i s   n o t   a   v a l i d   t i m e s t a m p  ' % s '   i s   n o t   a   v a l i d   G U I D   v a l u e  I n v a l i d   a r g u m e n t   t o   d a t e   e n c o d e  O u t   o f   m e m o r y  I / O   e r r o r   % d  T o o   m a n y   o p e n   f i l e s  F i l e   a c c e s s   d e n i e d  R e a d   b e y o n d   e n d   o f   f i l e 	 D i s k   f u l l  D u p l i c a t e s   n o t   a l l o w e d , S p e c i f i e d   L o g i n   C r e d e n t i a l   S e r v i c e   n o t   f o u n d " % s   ( V e r s i o n   % d . % d ,   B u i l d   % d ,   % 5 : s ) : % s   S e r v i c e   P a c k   % 4 : d   ( V e r s i o n   % 1 : d . % 2 : d ,   B u i l d   % 3 : d ,   % 5 : s )  3 2 - b i t   E d i t i o n  6 4 - b i t   E d i t i o n  W i n d o w s  W i n d o w s   V i s t a  W i n d o w s   S e r v e r   2 0 0 8 	 W i n d o w s   7  W i n d o w s   S e r v e r   2 0 0 8   R 2  W i n d o w s   2 0 0 0 
 W i n d o w s   X P  W i n d o w s   S e r v e r   2 0 0 3  W i n d o w s   S e r v e r   2 0 0 3   R 2  O b s e r v e r   i s   n o t   s u p p o r t e d  I n v a l i d   T i m e s p a n   f o r m a t  T i m e s p a n   e l e m e n t   t o o   l o n g  ' % s '   � r   i n g e t   g i l t i g t   d a t u m # ' % s '   � r   i n g e t   g i l t i g t   d a t u m   o c h   t i d # ' ' % s ' '   i s   n o t   a   v a l i d   i n t e g e r   v a l u e  ' % s '   � r   i n g e n   g i l t i g   t i d  I n v a l i d   a r g u m e n t   t o   t i m e   e n c o d e # N o   c o n t e x t - s e n s i t i v e   h e l p   i n s t a l l e d  N o   h e l p   f o u n d   f o r   c o n t e x t   % d  U n a b l e   t o   o p e n   I n d e x  U n a b l e   t o   o p e n   S e a r c h " U n a b l e   t o   f i n d   a   T a b l e   o f   C o n t e n t s $ N o   t o p i c - b a s e d   h e l p   s y s t e m   i n s t a l l e d  N o   h e l p   f o u n d   f o r   % s  A r g u m e n t   o u t   o f   r a n g e  I t e m   n o t   f o u n d     T h e   s p e c i f i e d   p a t h   w a s   n o t   f o u n d   T h e   p a t h   f o r m a t   i s   n o t   s u p p o r t e d  T h e   d r i v e   c a n n o t   b e   f o u n d   T h e   s p e c i f i e d   f i l e   w a s   n o t   f o u n d W T h e   g i v e n   " % s "   l o c a l   t i m e   i s   i n v a l i d   ( s i t u a t e d   w i t h i n   t h e   m i s s i n g   p e r i o d   p r i o r   t o   D S T ) . $ N o   h e l p   v i e w e r   t h a t   s u p p o r t s   f i l t e r s 7 S t r i n g   i n d e x   o u t   o f   r a n g e   ( % d ) .     M u s t   b e   > =   1   a n d   < =   % d \ I n v a l i d   U T F 3 2   c h a r a c t e r   v a l u e .     M u s t   b e   > =   0   a n d   < =   $ 1 0 F F F F ,   e x c l u d i n g   s u r r o g a t e   p a i r   r a n g e s r H i g h   s u r r o g a t e   c h a r   w i t h o u t   a   f o l l o w i n g   l o w   s u r r o g a t e   c h a r   a t   i n d e x :   % d .   C h e c k   t h a t   t h e   s t r i n g   i s   e n c o d e d   p r o p e r l y r L o w   s u r r o g a t e   c h a r   w i t h o u t   a   p r e c e d i n g   h i g h   s u r r o g a t e   c h a r   a t   i n d e x :   % d .   C h e c k   t h a t   t h e   s t r i n g   i s   e n c o d e d   p r o p e r l y 2 L e n g t h   o f   S t r i n g s   a n d   O b j e c t s   a r r a y s   m u s t   b e   e q u a l  I n v a l i d   T i m e o u t   v a l u e :   % s  T i m e s p a n   t o o   l o n g b T h e   d u r a t i o n   c a n n o t   b e   r e t u r n e d   b e c a u s e   t h e   a b s o l u t e   v a l u e   e x c e e d s   t h e   v a l u e   o f   T T i m e S p a n . M a x V a l u e  V a l u e   c a n n o t   b e   N a N 3 N e g a t i n g   t h e   m i n i m u m   v a l u e   o f   a   T i m e s p a n   i s   i n v a l i d    S t r i n g   e x p e c t e d  % s   e x p e c t e d $ % s   n o t   i n   a   c l a s s   r e g i s t r a t i o n   g r o u p  P r o p e r t y   % s   d o e s   n o t   e x i s t  S t r e a m   w r i t e   e r r o r  T h r e a d   c r e a t i o n   e r r o r :   % s  T h r e a d   E r r o r :   % s   ( % d ) - C a n n o t   t e r m i n a t e   a n   e x t e r n a l l y   c r e a t e d   t h r e a d , C a n n o t   w a i t   f o r   a n   e x t e r n a l l y   c r e a t e d   t h r e a d 2 C a n n o t   c a l l   S t a r t   o n   a   r u n n i n g   o r   s u s p e n d e d   t h r e a d ; C a n n o t   c a l l   C h e c k T e r m i n a t e d   o n   a n   e x t e r n a l l y   c r e a t e d   t h r e a d 9 C a n n o t   c a l l   S e t R e t u r n V a l u e   o n   a n   e x t e r n a l l y   c r e a t e   t h r e a d ' P a r a m e t e r   % s   c a n n o t   b e   a   n e g a t i v e   v a l u e * I n p u t   b u f f e r   e x c e e d e d   f o r   % s   =   % d ,   % s   =   % d  I n v a l i d   c h a r a c t e r s   i n   p a t h  T h e   s p e c i f i e d   p a t h   i s   t o o   l o n g  L i s t   i n d e x   o u t   o f   b o u n d s   ( % d ) + O u t   o f   m e m o r y   w h i l e   e x p a n d i n g   m e m o r y   s t r e a m ) % s   h a s   n o t   b e e n   r e g i s t e r e d   a s   a   C O M   c l a s s  N u m b e r   e x p e c t e d  A N S I   o r   U T F 8   e n c o d i n g   e x p e c t e d  % s   o n   l i n e   % d  E r r o r   r e a d i n g   % s % s % s :   % s  S t r e a m   r e a d   e r r o r  P r o p e r t y   i s   r e a d - o n l y  F a i l e d   t o   c r e a t e   k e y   % s  F a i l e d   t o   g e t   d a t a   f o r   ' % s '  I n v a l i d   c o m p o n e n t   r e g i s t r a t i o n  F a i l e d   t o   s e t   d a t a   f o r   ' % s '  R e s o u r c e   % s   n o t   f o u n d  % s . S e e k   n o t   i m p l e m e n t e d $ O p e r a t i o n   n o t   a l l o w e d   o n   s o r t e d   l i s t  C a n n o t   o p e n   f i l e   " % s " .   % s  I d e n t i f i e r   e x p e c t e d  U n a b l e   t o   w r i t e   t o   % s  I n v a l i d   b i n a r y   v a l u e  I n v a l i d   f i l e   n a m e   -   % s  I n v a l i d   s t r e a m   f o r m a t  ' % s '   i s   a n   i n v a l i d   m a s k   a t   ( % d ) $ ' ' % s ' '   i s   n o t   a   v a l i d   c o m p o n e n t   n a m e  I n v a l i d   p r o p e r t y   v a l u e  I n v a l i d   p r o p e r t y   p a t h  I n v a l i d   p r o p e r t y   v a l u e  I n v a l i d   d a t a   t y p e   f o r   ' % s '  I n v a l i d   s t r i n g   c o n s t a n t  L i n e   t o o   l o n g   L i s t   c a p a c i t y   o u t   o f   b o u n d s   ( % d )  L i s t   c o u n t   o u t   o f   b o u n d s   ( % d )    O L E   e r r o r   % . 8 x . M e t h o d   ' % s '   n o t   s u p p o r t e d   b y   a u t o m a t i o n   o b j e c t / V a r i a n t   d o e s   n o t   r e f e r e n c e   a n   a u t o m a t i o n   o b j e c t 7 D i s p a t c h   m e t h o d s   d o   n o t   s u p p o r t   m o r e   t h a n   6 4   p a r a m e t e r s  A n c e s t o r   f o r   ' % s '   n o t   f o u n d  C a n n o t   a s s i g n   a   % s   t o   a   % s  B i t s   i n d e x   o u t   o f   r a n g e * C a n ' t   w r i t e   t o   a   r e a d - o n l y   r e s o u r c e   s t r e a m  ' ' % s ' '   e x p e c t e d E C h e c k S y n c h r o n i z e   c a l l e d   f r o m   t h r e a d   $ % x ,   w h i c h   i s   N O T   t h e   m a i n   t h r e a d  C l a s s   % s   n o t   f o u n d  A   c l a s s   n a m e d   % s   a l r e a d y   e x i s t s % L i s t   d o e s   n o t   a l l o w   d u p l i c a t e s   ( $ 0 % x ) # A   c o m p o n e n t   n a m e d   % s   a l r e a d y   e x i s t s % S t r i n g   l i s t   d o e s   n o t   a l l o w   d u p l i c a t e s  C a n n o t   c r e a t e   f i l e   " % s " .   % s    I n v a l i d   i n d e x  U n a b l e   t o   i n s e r t   a n   i t e m  I n v a l i d   o w n e r  R i c h E d i t   l i n e   i n s e r t i o n   e r r o r  F a i l e d   t o   L o a d   S t r e a m  F a i l e d   t o   S a v e   S t r e a m   % s   i s   a l r e a d y   a s s o c i a t e d   w i t h   % s E % d   i s   a n   i n v a l i d   P a g e I n d e x   v a l u e .     P a g e I n d e x   m u s t   b e   b e t w e e n   0   a n d   % d = T h i s   c o n t r o l   r e q u i r e s   v e r s i o n   4 . 7 0   o r   g r e a t e r   o f   C O M C T L 3 2 . D L L  D a t e   e x c e e d s   m a x i m u m   o f   % s  D a t e   i s   l e s s   t h a n   m i n i m u m   o f   % s 4 Y o u   m u s t   b e   i n   S h o w C h e c k b o x   m o d e   t o   s e t   t o   t h i s   d a t e # F a i l e d   t o   s e t   c a l e n d a r   d a t e   o r   t i m e % F a i l e d   t o   s e t   m a x i m u m   s e l e c t i o n   r a n g e $ F a i l e d   t o   s e t   c a l e n d a r   m i n / m a x   r a n g e % F a i l e d   t o   s e t   c a l e n d a r   s e l e c t e d   r a n g e    I n v a l i d   s t y l e   h a n d l e  I n v a l i d   s t y l e   f o r m a t  V C L   S t y l e   F i l e % C l a s s   ' % s '   i s   n o t   r e g i s t e r e d   f o r   ' % s '  % s   p a r a m e t e r   c a n n o t   b e   n i l 0 A   S t y l e H o o k   c l a s s   h a s   n o t   b e e n   r e g i s t e r e d   f o r   % s # F e a t u r e   n o t   s u p p o r t e d   b y   t h i s   s t y l e  F a i l e d   t o   c l e a r   t a b   c o n t r o l   F a i l e d   t o   d e l e t e   t a b   a t   i n d e x   % d " F a i l e d   t o   r e t r i e v e   t a b   a t   i n d e x   % d   F a i l e d   t o   g e t   o b j e c t   a t   i n d e x   % d " F a i l e d   t o   s e t   t a b   " % s "   a t   i n d e x   % d   F a i l e d   t o   s e t   o b j e c t   a t   i n d e x   % d < M u l t i L i n e   m u s t   b e   T r u e   w h e n   T a b P o s i t i o n   i s   t p L e f t   o r   t p R i g h t  I n v a l i d   i t e m   l e v e l   a s s i g n m e n t   I n v a l i d   l e v e l   ( % d )   f o r   i t e m   " % s "  U T F - 7 % C a n n o t   r e m o v e   s h e l l   n o t i f i c a t i o n   i c o n " P a g e C o n t r o l   m u s t   f i r s t   b e   a s s i g n e d " % s   r e q u i r e s   W i n d o w s   V i s t a   o r   l a t e r  B u t t o n % d  R a d i o B u t t o n % d  C a p t i o n   c a n n o t   b e   e m p t y : C a t e g o r y P a n e l   m u s t   h a v e   a   C a t e g o r y P a n e l G r o u p   a s   i t s   p a r e n t = O n l y   C a t e g o r y P a n e l s   c a n   b e   i n s e r t e d   i n t o   a   C a t e g o r y P a n e l G r o u p  N o   h e l p   k e y w o r d   s p e c i f i e d .  U n a b l e   t o   l o a d   s t y l e   ' % s '  U n a b l e   t o   l o a d   s t y l e s :   % s  S t y l e   ' % s '   a l r e a d y   r e g i s t e r e d # S t y l e   c l a s s   ' % s '   a l r e a d y   r e g i s t e r e d  S t y l e   ' % s '   n o t   f o u n d  S t y l e   c l a s s   ' % s '   n o t   f o u n d   7 L e n g t h   o f   v a l u e   a r r a y   m u s t   b e   > =   l e n g t h   o f   p r o m p t   a r r a y  P r o m p t   a r r a y   m u s t   n o t   b e   e m p t y 	 & U s e r n a m e 	 & P a s s w o r d  & D o m a i n  L o g i n 	 S e p a r a t o r  E r r o r   s e t t i n g   % s . C o u n t 8 L i s t b o x   ( % s )   s t y l e   m u s t   b e   v i r t u a l   i n   o r d e r   t o   s e t   C o u n t # N o   O n G e t I t e m   e v e n t   h a n d l e r   a s s i g n e d  " % s "   i s   a n   i n v a l i d   p a t h  A N S I  A S C I I  U n i c o d e  B i g   E n d i a n   U n i c o d e  U T F - 8     C l i p b o a r d   d o e s   n o t   s u p p o r t   I c o n s  C a n n o t   o p e n   c l i p b o a r d :   % s  T e x t   e x c e e d s   m e m o   c a p a c i t y + O p e r a t i o n   n o t   s u p p o r t e d   o n   s e l e c t e d   p r i n t e r . T h e r e   i s   n o   d e f a u l t   p r i n t e r   c u r r e n t l y   s e l e c t e d / M e n u   ' % s '   i s   a l r e a d y   b e i n g   u s e d   b y   a n o t h e r   f o r m  P i c t u r e :    ( % d x % d )  P r e v i e w  C a n n o t   o p e n   A V I  D o c k e d   c o n t r o l   m u s t   h a v e   a   n a m e % E r r o r   r e m o v i n g   c o n t r o l   f r o m   d o c k   t r e e    -   D o c k   z o n e   n o t   f o u n d    -   D o c k   z o n e   h a s   n o   c o n t r o l L E r r o r   l o a d i n g   d o c k   z o n e   f r o m   t h e   s t r e a m .   E x p e c t i n g   v e r s i o n   % d ,   b u t   f o u n d   % d . , M u l t i s e l e c t   m o d e   m u s t   b e   o n   f o r   t h i s   f e a t u r e  E n d  H o m e  L e f t  U p  R i g h t  D o w n  I n s  D e l  S h i f t +  C t r l +  A l t +  ( N o n e )  V a l u e   m u s t   b e   b e t w e e n   % d   a n d   % d  A l l  U n a b l e   t o   i n s e r t   a   l i n e  I n v a l i d   c l i p b o a r d   f o r m a t  A v b r y t  & H j � l p  & A v b r y t  & F � r s � k   i g e n 	 & I g n o r e r a  & A l l a  N & e j   t i l l   a l l a  J & a   t i l l   a l l a  & S t � n g  B k S p  T a b  E s c  E n t e r  S p a c e  P g U p  P g D n  T I F F   I m a g e s  G r i d   t o o   l a r g e   f o r   o p e r a t i o n   T o o   m a n y   r o w s   o r   c o l u m n s   d e l e t e d  G r i d   i n d e x   o u t   o f   r a n g e 1 F i x e d   c o l u m n   c o u n t   m u s t   b e   l e s s   t h a n   c o l u m n   c o u n t + F i x e d   r o w   c o u n t   m u s t   b e   l e s s   t h a n   r o w   c o u n t & C a n n o t   i n s e r t   o r   d e l e t e   r o w s   f r o m   g r i d  O g i l t i g t   i n p u t v � r d e 9 O g i l t i g t   i n p u t v � r d e .   A n v � n d   E S C   f � r   a t t   a v b r y t a   � n d r i n g a r  V a r n i n g  F e l  I n f o r m a t i o n  B e k r � f t a  & J a  & N e j  O K  & N o  & H e l p  & C l o s e  & I g n o r e  & R e t r y  A b o r t  & A l l  C a n n o t   d r a g   a   f o r m " A n   e r r o r   r e t u r n e d   f r o m   D D E     ( $ 0 % x ) / D D E   E r r o r   -   c o n v e r s a t i o n   n o t   e s t a b l i s h e d   ( $ 0 % x ) 0 E r r o r   o c c u r r e d   w h e n   D D E   r a n   o u t   o f   m e m o r y   ( $ 0 % x ) " U n a b l e   t o   c o n n e c t   D D E   c o n v e r s a t i o n 	 M e t a f i l e s  E n h a n c e d   M e t a f i l e s  I c o n s  B i t m a p s  M e n u   i n d e x   o u t   o f   r a n g e  M e n u   i n s e r t e d   t w i c e  S u b - m e n u   i s   n o t   i n   m e n u  N o t   e n o u g h   t i m e r s   a v a i l a b l e ! P r i n t e r   i s   n o t   c u r r e n t l y   p r i n t i n g  P r i n t i n g   i n   p r o g r e s s  P r i n t e r   i n d e x   o u t   o f   r a n g e  P r i n t e r   s e l e c t e d   i s   n o t   v a l i d  % s   o n   % s @ G r o u p I n d e x   c a n n o t   b e   l e s s   t h a n   a   p r e v i o u s   m e n u   i t e m ' s   G r o u p I n d e x 5 C a n n o t   c r e a t e   f o r m .   N o   M D I   f o r m s   a r e   c u r r e n t l y   a c t i v e 0 C a n   o n l y   m o d i f y   a n   i m a g e   i f   i t   c o n t a i n s   a   b i t m a p * A   c o n t r o l   c a n n o t   h a v e   i t s e l f   a s   i t s   p a r e n t  O K  A v b r y t  & Y e s    I n v a l i d   i m a g e   s i z e  I n v a l i d   I m a g e L i s t  U n a b l e   t o   R e p l a c e   I m a g e  I n v a l i d   I m a g e L i s t   I n d e x ) F a i l e d   t o   r e a d   I m a g e L i s t   d a t a   f r o m   s t r e a m ( F a i l e d   t o   w r i t e   I m a g e L i s t   d a t a   t o   s t r e a m $ E r r o r   c r e a t i n g   w i n d o w   d e v i c e   c o n t e x t  E r r o r   c r e a t i n g   w i n d o w   c l a s s + C a n n o t   f o c u s   a   d i s a b l e d   o r   i n v i s i b l e   w i n d o w ! C o n t r o l   ' % s '   h a s   n o   p a r e n t   w i n d o w $ P a r e n t   g i v e n   i s   n o t   a   p a r e n t   o f   ' % s '  C a n n o t   h i d e   a n   M D I   C h i l d   F o r m ) C a n n o t   c h a n g e   V i s i b l e   i n   O n S h o w   o r   O n H i d e " C a n n o t   m a k e   a   v i s i b l e   w i n d o w   m o d a l  S c r o l l b a r   p r o p e r t y   o u t   o f   r a n g e  % s   p r o p e r t y   o u t   o f   r a n g e 0 T a b   p o s i t i o n   i n c o m p a t i b l e   w i t h   c u r r e n t   t a b   s t y l e 0 T a b   s t y l e   i n c o m p a t i b l e   w i t h   c u r r e n t   t a b   p o s i t i o n  B i t m a p   i m a g e   i s   n o t   v a l i d  I c o n   i m a g e   i s   n o t   v a l i d  M e t a f i l e   i s   n o t   v a l i d  I n v a l i d   p i x e l   f o r m a t  I n v a l i d   i m a g e  S c a n   l i n e   i n d e x   o u t   o f   r a n g e ! C a n n o t   c h a n g e   t h e   s i z e   o f   a n   i c o n % C a n n o t   c h a n g e   t h e   s i z e   o f   a   W I C   I m a g e   I n v a l i d   o p e r a t i o n   o n   T O l e G r a p h i c $ U n k n o w n   p i c t u r e   f i l e   e x t e n s i o n   ( . % s )  U n s u p p o r t e d   c l i p b o a r d   f o r m a t  O u t   o f   s y s t e m   r e s o u r c e s  C a n v a s   d o e s   n o t   a l l o w   d r a w i n g # T e x t   f o r m a t   f l a g   ' % s '   n o t   s u p p o r t e d   ��ߘ{<:y&q?	*%TPF0TAboutDialogAboutDialogLeftuTop{HelpType	htKeywordHelpKeywordui_aboutBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption	Om WinSCPClientHeight�ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenter
DesignSize�� PixelsPerInch`
TextHeight TLabelApplicationLabelLeftHTopWidth4HeightCaptionApplication  TLabelVersionLabelLeftHTopWidthHeightCaptionVersion 2.0.0 (Build 12) XX  TLabelWinSCPCopyrightLabelLeftHTop8Width� HeightCaption%   Copyright © 2000-2003 Martin Prikryl  TLabelProductSpecificMessageLabelLeftHTopdWidthHeightCaption5   För att skicka in kommentarer och rapportera buggar:  TLabelTranslatorLabelLeftHTop� WidthJHeightCaptionTranslatorLabel  TImageImageLeftTopWidth1Height Center	Picture.Data
� TIcon         h  v        �	  �         �  f  **         00     �%  <  @@     (B  �a  ��     ( �  (                                     jjj�iii�iii�iii�iii�iii�jjj�E�E�T�T�^�_�i�i�s�t�~�~���������k�kXiii���������������������iii�2�4aE�E�����������-�-�����iii���������������������iii��D 2�4aD�E��� �� �� ��������iii���������������������iii��D 0�2;=�>�	�
� �� �� ����~�~�jjj�iii�iii�iii�iii�iii�jjj�� 7)�*��� �� �� �� ����s�t��D fff������D ����fff�]�[��	�� �� �� ��	�
�����i�i��u%	fff������D ����fff�]���� �� �� ����=�>�D�E���^�_��}8�fff�������������fff��z	�/�� �� ��	��(�*�-�.@5�7[E�F�T�T��A��sg�fff�fff�fff�q^��o ��v �-�������<�D �D 5�7[D�E��G��a��}9��5��l��f ��j ��o ��{	�Z��X�^�D �D �D �D 2�3�M��R��X��^	��] ��a ��f ��r����9�D �D �D �D �D �D �R��M��O ��S ��X ��] ��l��*��}!:�D �D �D �D �D �D �D ��X��I��J ��O ��S ��^	��5��}-:�D �D �D �D �D �D �D �D �^��E��E ��J ��O ��X��}9��}2T�D �D �D �D �D �D �D �D �~[��X%��E��I��M��R��a��~:��{0S�D �D �D �D �D �D �D �rOO�~[��^���X��R��M��G��A��}8��u%	�D �D �D �D �D �D       �  �     �   �          ?      �  �  �   �  �  (      0                              ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �Հo�suR�V�M�Q�L�P�L�P�K�P�L�Q�Y�`�'=':   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���b�f��� � � � � � � � � � �� �m�r�   ��� ��� ��� ���                               ^�a��� � � � � � ���>�>�m�r�   ��� ��� ��� ���    CCC"777A111I111I444I444I777J777J777J999LRlTa>�A� � � � ���4�4�>�>�n�q�   ��� ��� ��� ��� ��� ttt�\\\�ggg�fff�mmm�www�zzz�yyy�}}}�����V�X��� � ���*�*�3�3�=�=�m�q�   ��� ��� ��� ��� ���+DDD�(((�222�???�???�===�EEE�CCC�KMK�I}J� �!�������)�)�3�3�<�<�n�q�   ��� ��� ��� ��� ���+JJJ�,,,�777�GGG�HHH�EEE�PPP�MMM�I]I�?u@�6�7�'�(�'�(�!�"�C�D�;�;�<�<�n�q�   ��� ��� ��� ��� ���*GGG�333�>>>�NNN�QQQ�MMM�\\\�VVV�Y]Y�VsW�Q�R�B�C�:�;�L�N�k�nfv�x�D�D�p�s�   
��� ��� ��� ��� ���)AAA�999�DDD�TTT�YYY�SSS�fff�___�ddd�ptp�o�p�Z�[�\�]�����   ���z�}�}び   ��� ��� ��� ��� ���)KKK�@@@�III�ZZZ�```�XXX�ppp�hhh�kkk�}}}�����w�x�x�y�����   ��� ��������� ��� ��� ��� ��� ���(OOO�GGG�MMM�___�ccc�]]]�zzz�qqq�sss�������������xxx�����   ��� ��� ��� ��� ��� ��� ��� ��� ���&PPP�MMM�RRR�bbb�eee�aaa�����xxx�|||���������������������   ��� ��� ��� ���          ��� ���ZZZ�TTT�VVV�eee�ggg�fff�����������������������������v   ��� ��� ��� ��� udW0)$      ������w���򦦦��������Ͷ��������������ƭ������������������"   ��� ��� ��� ��� �uf�f�   �|b��CrwlZ���������GD<Y            	��������eee�      ��� ��� ��� ��� ��� ��R��q��a�r\I:�F��} �|mW���������lX0jRF+   ���    	��������eee�      ��� ��� ��� ��� ��� �L��i ��p��@��v ��x ��mU����������n;��oO         ��������eee�      ��� ��� ��� ��� ��� �G��d ��i ��m ��r ��xËnO���������qj`�   '      /�����ccc�      ��� ��� ��� ��� ��� �C��` ��d ��i ��r��x
��}1թ�����������kkk�jjj�jjj�qqq򨨨�����^^^�   ��� ��� ��� ��� ��� ��� �}>��[ ��` ��j
��q��s
��4؎�������������������������������ggg�      ��� ��� ��� ��� ��� ��� �y;��V ��d��l��m��o
��t��s�zzyā��쒒�򅅅�ttt�lll�eee�+++   ��� ��� ��� ��� ��� ��� ��� ށJr�_��f��h��j��k��m��r��f�(!   	               ��� ��� ��� ��� ��� ��� ��� ��� ��cބN��D���B��B��B��B���C���b�䵔   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �� �� �� �� �  �  �  �  �  �  �  �  � ? � ? �| |  <  <      �  � �� �� (       @                              ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���          
                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    +t�{Ql�qhg�nme�loc�jqa�gt_�ev\�ct/A   *      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��>h�l�*�,�"�$�"�$�"�$�"�$�"�$�"�%�$�&�Q�V�i�p�   (   ��� ��� ��� ��� ��� ��� ��� ���                               f�fw�|��� � � � � � � � � � � � � � ���m�p�@lFP   ��� ��� ��� ��� ��� ���             	   	   	   	   	   	   	   	   	   	(;(t�y��� � � � � � � � � � ���=�=�I�I�{ނ�   ��� ��� ��� ��� ���             !   %   &   &   &   &   &   &   &   &   &   &+q�t��� � � � � � ���5�5�<�<�D�D�~ᄺ   ��� ��� ��� ��� ���    rrr���^vvv�zzz�vvv�vvv�zzz������������������������������O�Q� � � � � � ���-�-�5�5�<�<�D�D�ⅸ   ��� ��� ��� ��� ���    ���rTTT�FFF�PPP�RRR�PPP�VVV�___�eee�ggg�fff�jjj�ooo�w}w�U�W��� � � � ���&�&�-�-�4�4�<�<�C�C��ᄷ   ��� ��� ��� ��� ���    ����111�&&&�000�666�>>>�===�;;;�???�DDD�BBB�FFF�QUQ�J�K� �!���	�
�	�	���&�&�-�-�4�4�;�;�C�C��ᅶ   ��� ��� ��� ��� ���    ����444�'''�333�:::�FFF�EEE�AAA�FFF�MMM�JJJ�KLK�HkI�6x7�/�0�"�#���!�"���%�%�,�,�4�4�;�;�B�B��↵   ��� ��� ��� ��� ���    ����777�+++�999�>>>�KKK�MMM�GGG�NNN�UUU�PPP�OWO�IfJ�GwH�A�B�5�6�1�2�.�/�)�*�9�9����B�C�;�;�B�B��㈲   ��� ��� ��� ��� ���    ����555�000�@@@�CCC�QQQ�TTT�LLL�SSS�]]]�XXX�YYY�[f[�Zw[�V�W�I�J�?�@�=�>�J�L�v�x�;O;�副I�J�C�C��犪   ��� ��� ��� ��� ���    zzz�111�444�FFF�FFF�VVV�ZZZ�PPP�ZZZ�ddd�^^^�___�ggg�nyn�n�o�\�]�N�O�V�W��à�      ����䋱s�t��މ?   ��� ��� ��� ��� ���    ����666�888�KKK�JJJ�ZZZ�___�UUU�___�lll�eee�fff�mmm�}}}�����r�s�d�e�������      ��� �����      ��� ��� ��� ��� ���    ����<<<�===�QQQ�MMM�^^^�ccc�XXX�eee�ttt�jjj�lll�rrr�����������������vvv�����      ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ����<<<�@@@�XXX�OOO�aaa�eee�\\\�jjj�{{{�qqq�rrr�www�����������������www�����      ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ����===�EEE�^^^�PPP�ccc�ggg�^^^�nnn�����www�xxx�~~~�������������������������      ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ����>>>�KKK�ddd�RRR�fff�jjj�___�sss�����|||�|||�����������������������������      ��� ��� ��� ��� ���             ���    ���dfff�bbb�{{{�eee�xxx�{{{�ppp�������������}}}����������������������������y      ��� ��� ��� ��� ���    �vh            ������r���У���������������������č��ʈ�����������ŷ������������������s���"   ��� ��� ��� ��� ��� ��� ��}���͞~eD         ��t(�Ju�t?���������~~~�KICp               cccq��������xxx�R      ��� ��� ��� ��� ��� ��� ��� ��~��s��[͑u^K   ��j8�N�� ��u;���������~~~�`U<z6)	      ���    cccq��������xxx�Q      ��� ��� ��� ��� ��� ��� ��� ��m��k ��m ��Zͽ�yq�O��z ��{ ��v7���������~~~�r^7��k0|sa
   ���    cccq��������xxx�Q      ��� ��� ��� ��� ��� ��� ��� �h��f ��j ��m ���/��s ��w ��x ��w5���������~~~��k=���\:            aaat��������xxx�   O      ��� ��� ��� ��� ��� ��� ��� �c��c ��f ��j ��m ��q ��s ��y��w,Ƭ�����������~te�   -            ^^^���������vvv�A      ��� ��� ��� ��� ��� ��� ��� �^��` ��c ��f ��j ��m ��u��x	��}�����������vvv�[[[�RRR�SSS�SSS�WWW�eee���������lll�   ,      ��� ��� ��� ��� ��� ��� ��� �Z��\ ��` ��c ��f ��o	��t��v	��Ѝ�}���������������������������������������������ddd�         ��� ��� ��� ��� ��� ��� ��� �U��Y ��\ ��` ��j��o��q��r	���"�հ������������������������������������������ggg�+++0      ��� ��� ��� ��� ��� ��� ��� ��� �Q��U ��Y ��e��l��m��n��p	��t��nԤ��{���蒒��������������xxx�uuu�mmm�eee�+++$   	   ��� ��� ��� ��� ��� ��� ��� ��� ��� �Xw�Z��`��h��i��j��k��l
��n��t	���jӴ��VZZZ            	      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ́[
�O��g��e��f��g��i��i
��j��m��o ���m�׭�5                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �f�Z��O��P��Q��S��U��V���W���a����o��|
   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���������������������  �  �  �  �  �  !�  s�  {�  �  �  �  �  �� �������� �� ��  �  �  �  ����������(   *   T                              ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                       ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                   "   $   &   (   *   ,   .   /   ,   $         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       �ܑ:�ꇶ}��|��{��{��z��z��z��y��y��{��s�|�5T8R   ,      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���xg�j��� � � � � � � � � � � � � � � � � � � � ������HtN\   "   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                     ����茯#�$� � � � � � � � � � � � � � � � � � � � ���J�K����   )   ��� ��� ��� ��� ��� ��� ��� ��� ���                                                 V�V�拰!�#� � � � � � � � � � � � � � � � ���=�=�C�C�����-   ��� ��� ��� ��� ��� ��� ���                                                          &:&�ሴ �"� � � � � � � � � � � � ���7�7�=�=�C�C�����*1   ��� ��� ��� ��� ��� ��� ���       	      #   ,   /   0   0   0   0   0   0   0   0   0   0   0   0   0   1:���	�	� � � � � � � � ���1�1�7�7�=�=�B�B����+0   ��� ��� ��� ��� ��� ���       DDD���Fuuu^jjjjhhhnhhhnjjjolllolllommmpmmmpoooqppprppprrrrrssssssssuuutwwwv�Ê�.�0� � � � � � � � ���,�,�2�2�7�7�=�=�B�B����-.   ��� ��� ��� ��� ��� ���       ���Mttt�]]]�ccc�mmm�mmm�hhh�^^^�ppp��������������������������������������;�<��� � � � � � ���&�&�,�,�1�1�7�7�<�<�B�B����/,   ��� ��� ��� ��� ��� ���       ����GGG��***�111�444�===�>>>�<<<�888�888�???�@@@�>>>�AAA�DDD�IJI�e{e�8�9������� � �
�
� � �&�&�,�,�1�1�6�6�<�<�B�B����1*   ��� ��� ��� ��� ��� ���       ����HHH��)))�000�333�===�AAA�@@@�<<<�===�EEE�FFF�DDD�FFF�JJJ�Zh[�=�>�&�'����������� � �&�&�+�+�1�1�6�6�<�<�A�A���� 3 (   ��� ��� ��� ��� ��� ���       ����LLL��+++�444�777�AAA�HHH�EEE�AAA�AAA�KKK�LLL�JJJ�KKK�PWP�BoC�6v7�2�3�+�,�� ���� � �!� � �%�%�+�+�0�0�6�6�<�<�A�A����"6"&   ��� ��� ��� ��� ��� ���       ����SSS�   �000�888�999�EEE�NNN�KKK�EEE�FFF�RRR�SSS�OOO�OQO�I^I�EiF�CuD�@�A�8�9�-�.�-�.�(�)�.�/�"�#�'�'�{�~�K�L�6�6�;�;�A�A����$:$#   ��� ��� ��� ��� ��� ���       ����NNN�"""�444�===�===�JJJ�RRR�PPP�III�JJJ�WWW�YYY�UUU�TTT�T\T�RhR�QuR�O�P�G�H�?�@�9�:�1�2�<�=�-�.�u�wۄƈB�银O�P�;�;�@�@����-H-   	��� ��� ��� ��� ��� ���       ����FFF�$$$�888�BBB�@@@�NNN�VVV�VVV�MMM�NNN�]]]�___�ZZZ�ZZZ�]]]�_g_�^t^�_�`�Y�Z�M�N�E�F�<�=�J�K�{�}�d�hE   V�V	�엶T�U�@�@���� 0    ��� ��� ��� ��� ��� ���       ����???�&&&�<<<�GGG�CCC�QQQ�ZZZ�ZZZ�PPP�QQQ�ccc�fff�___�___�bbb�hhh�nvn�q�q�j�k�Z�[�Q�R�G�H���������       	   ����혷a�c���      ��� ��� ��� ��� ��� ���       ����HHH�'''�@@@�KKK�DDD�TTT�]]]�___�TTT�UUU�iii�kkk�ccc�eee�eee�mmm�yyy�����~�~�i�j�`�a�o�p��������r      	   ��� �ے�񞽙�9   ��� ��� ��� ��� ��� ��� ���       ����QQQ�)))�EEE�PPP�FFF�WWW�aaa�aaa�WWW�WWW�nnn�qqq�iii�iii�jjj�qqq����������y�y�z�z�xzx��������q      	   ��� ��� ������ ��� ��� ��� ��� ��� ��� ��� ���       ����UUU�+++�HHH�TTT�GGG�YYY�ddd�ddd�YYY�ZZZ�ttt�www�nnn�nnn�ooo�vvv���������������������xxx��������q      	   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ����UUU�---�MMM�YYY�III�[[[�fff�eee�\\\�\\\�yyy�|||�rrr�sss�uuu�yyy���������������������zzz��������p      	   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ����WWW�...�PPP�```�KKK�^^^�iii�ggg�^^^�___�~~~�����vvv�vvv�xxx�}}}���������������������}}}��������n         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ����WWW�000�UUU�eee�LLL�___�jjj�ggg�^^^�aaa���������zzz�{{{�}}}�����������������������������󙙙i         ��� ��� ��� ��� ��� ��� ���          ��� ��� ���    ���zYYY�222�YYY�jjj�KKK�```�kkk�iii�]]]�bbb���������������������������������������|||�����\         ��� ��� ��� ��� ��� ���                   ���    ���>zzz�ZZZ�zzz�����jjj�}}}���������yyy�����������������rrr������������������������������������Ϳ��C   	   ��� ��� ��� ��� ��� ��� ���    +% 
                  ������D��������������������������������ǔ��Ώ��̏���������������ܺ��������������������������K���      ��� ��� ��� ��� ��� ��� ���    ����Ϥ�^         	         
ֲ�P֒)ovn_Բ�����������fee�   7      
               	eee�������������hhh�   C   "      ��� ��� ��� ��� ��� ��� ��� ��� ��� �{j��n���Yռ�ui            ߶�c�.��} uyn]ش�����������ffe�0! @      	      ���       eee�������������hhh�   B       	   ��� ��� ��� ��� ��� ��� ��� ��� ��� �g��)��o ���Yظ�sm   "   ޲�z�0��~ ��{ �|o\۵�����������ffe�W; LQ8 &('$   ��� ���       eee�������������hhh�   B       	   ��� ��� ��� ��� ��� ��� ��� ��� ��� �z�y��l ��n ��Yٵ�qoګ���1��z ��{ ��z �~oZ߷�����������ffe�tL X�Y3��h   ��� ���       eee�������������hhh�   A       	   ��� ��� ��� ��� ��� ��� ��� ��� ��� 變z�u��i ��k ��n ���Y��2��u ��w ��y ��y ��oY㹹����������ffe��Zd��TMnfY               eee�������������hhh�   A      	   ��� ��� ��� ��� ��� ��� ��� ��� ��� �{z�r��f ��i ��k ��n ��p ��s ��u ��w ��y��pX溺����������hgf���N�KC:1         	   	      ccc�������������hhh�   =         ��� ��� ��� ��� ��� ��� ��� ��� ��� �wz�p��c ��f ��i ��k ��n ��p ��s ��x��z��tQⰰ����������www�WSNw9   )   #   !   !   #   (bbbӗ�����������fff�   7         ��� ��� ��� ��� ��� ��� ��� ��� ��� �r{�m��a ��c ��f ��i ��k ��n ��t��y
��x�̀1͓���������������qqq�YYY�EEE�GGG�GGG�GGG�GGG�^^^�fff�������������ddd�   -      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �n{�j��^ ��a ��c ��f ��i ��p	��u��v
��z��ˀ~}���������������������www�vvv�vvv�vvv�vvv���������������������bbb�         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �j{�g��\ ��^ ��a ��c ��l
��r��r��t
��x��ֻ��諫������������������������������������������������������ccc�)         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �f{�d��Y ��\ ��^ ��i��n��o��p��q
��t���J�ܹ�����Ӧ�����������������������������������������������bbb�SSSe         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �bz�b��V ��Y ��e��k��l��m��n��o
��p��x���k�ή������|||񁁁�������������|||�rrr�ppp�jjj�eee�eee�!         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �e]�d��T ��`��h��j��j��k��k��l��n��p	��w���f�Ѭ��ddd1mmm&eee2kkk@iiiAeee?XXX=UUU<                  ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ތc�~C��]��f��f��g��h��h��i��j��k��l��n��r���]�߱�q                              ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �_}ۃK��e��d��e��f��g��g��h��h	��j��k��m���!���ز�(                  ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �bB�a��^��`��b��d��f��i���k���m���o���u����w�      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ������  ������  �����  �����  ���� �  ���� �  ���� �  ���� �  ���� �  ��   �  �    �  �    �  �    �  �    �  �    �  �   p�  �   x�  �   ��  �   ��  �   ��  �   ��  �   ��  �   ��  ��  ��  ��  ��  �� ��  �����  �����  � ���  � ���  � ���  � ��  � ���  �  ��  �  ��  �  ��  �  ��  �  ?��  �����  �����  � ����  �����  (   0   `                              ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���          
                   !   #   %   &   (   )   *   (   #            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ~˃9�ڈp|ׁ�x�~�v�|�u�z�s�{�s�z�q�x�p�w�o�v�n�u�n�u�[�aq&C   0         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���퓮e�i�;�=�1�3�1�3�1�4�1�4�1�4�1�4�1�4�1�4�1�4�1�4�3�6�Q�W����W�]s   /      	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���씯*�,� � � � � � � � � � � � � � � � � � � � � � � � � � �������9_@P   !   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                 ���
�따*�,� � � � � � � � � � � � � � � � � � � � � � ���@�@�d�e�~ۅ�   %   ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                          VyV�鑳*�,� � � � � � � � � � � � � � � � � � ���;�;�A�A�K�K����   &   ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                +=+�⎹+�,� � � � � � � � � � � � � � ���6�6�<�<�@�@�E�E�����   %   ��� ��� ��� ��� ��� ��� ��� ���                '   ,   .   /   /   /   /   /   /   /   /   /   /   /   /   /   /   /   0 9����� � � � � � � � � � ���1�1�6�6�;�;�@�@�E�E�����   $   ��� ��� ��� ��� ��� ��� ��� ���       @@@$YYYDLLLTGGGZEEE]GGG]GGG]GGG]III^III^III^KKK_KKK_KKK_MMM_MMM_MMM_PPP`PPP`PPP`OOOa���S�U� � � � � � � � � � ���,�,�1�1�6�6�;�;�@�@�E�E�����   #   ��� ��� ��� ��� ��� ��� ���       ���+����|||�}}}��������􊊊�����yyy��������򦦦𦦦響��﨨�響��שּׁ����Ǳ�]�_��� � � � � � � � ���'�'�,�,�1�1�6�6�;�;�@�@�D�D�����   !   ��� ��� ��� ��� ��� ��� ���       ���Lhhh�...�***�333�777�;;;�AAA�BBB�BBB�>>>�???�@@@�CCC�CCC�BBB�EEE�GGG�KKK�OOO�gwh�N�P���	�
��� � � � �
�
�"�"�'�'�,�,�1�1�6�6�:�:�?�?�D�D�����      ��� ��� ��� ��� ��� ��� ���       ���Paaa��###�---�111�444�<<<�>>>�>>>�:::�999�<<<�BBB�CCC�AAA�CCC�EEE�JJJ�]h]�K�M�� �����	�
�������"�"�'�'�,�,�1�1�5�5�:�:�?�?�D�D�����      ��� ��� ��� ��� ��� ��� ���       ���Ohhh��###�---�111�444�>>>�CCC�DDD�>>>�>>>�@@@�HHH�HHH�FFF�GGG�KKK�W\W�I~J�-{.�)�*�"�#�����������"�"�'�'�,�,�0�0�5�5�:�:�?�?�D�D����      ��� ��� ��� ��� ��� ��� ���       ���Nooo��$$$�111�555�888�BBB�HHH�JJJ�BBB�AAA�EEE�MMM�NNN�KKK�KKK�MPM�GiH�:p;�8z9�3�4�,�-�"�#���#�$�#�$� �!�!�!�&�&�,�,�0�0�5�5�:�:�?�?�D�D�����      ��� ��� ��� ��� ��� ��� ���       ���Nuuu��'''�555�888�;;;�EEE�LLL�OOO�EEE�FFF�III�SSS�TTT�PPP�PPP�LZL�HeI�EnF�CyD�?�@�8�9�/�0�/�0�*�+�,�-�*�+�"�#�/�/����S�S�5�5�:�:�>�>�C�C����      ��� ��� ��� ��� ��� ��� ���       ���Mooo��)))�999�<<<�>>>�III�QQQ�TTT�JJJ�III�MMM�XXX�YYY�TTT�TTT�UYU�RcR�PmQ�PyQ�M�N�F�G�?�@�9�:�2�3�6�7�6�7�/�0��هلĈ<�혺V�W�9�9�>�>�C�C����      	��� ��� ��� ��� ��� ��� ���       ���Lddd��,,,�===�???�AAA�LLL�TTT�YYY�LLL�LLL�QQQ�]]]�^^^�YYY�YYY�ZZZ�^b^�\m\�]z^�[�\�V�W�J�K�D�E�;�<�A�B�H�I�΄�h�l;   ^�u�Z�[�>�>�D�E�����      ��� ��� ��� ��� ��� ��� ���       ���LXXX��...�BBB�CCC�CCC�OOO�XXX�___�PPP�PPP�UUU�ccc�ccc�]]]�^^^�^^^�eee�hlh�j{j�k�l�d�e�V�W�P�Q�D�E�O�P��̗�|�~a      	   �ȏ	��^�_�W�X���      ��� ��� ��� ��� ��� ��� ���       ���K[[[��111�FFF�FFF�DDD�RRR�ZZZ�bbb�SSS�RRR�WWW�iii�hhh�aaa�bbb�bbb�iii�ooo�z~z�{�{�t�u�c�d�\�]�P�Q���������cccN      	      ���򞽘����B      ��� ��� ��� ��� ��� ��� ���       ���Jhhh��333�JJJ�JJJ�FFF�UUU�]]]�eee�VVV�UUU�[[[�mmm�nnn�eee�fff�fff�mmm�ttt�������������q�r�j�k�s�s���������cccN      	   ��� ��� �����Z      ��� ��� ��� ��� ��� ��� ��� ���       ���Isss�!!!�555�NNN�MMM�HHH�WWW�___�ggg�XXX�WWW�^^^�rrr�sss�jjj�kkk�kkk�qqq�www�������������������yyy�yyy�����```M      	   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ���Ivvv�!!!�888�SSS�PPP�JJJ�YYY�aaa�jjj�[[[�YYY�aaa�www�xxx�nnn�nnn�nnn�uuu�{{{���������������������xxx�qqq�����```M      	   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ���Hvvv�"""�:::�XXX�TTT�KKK�[[[�ddd�lll�[[[�\\\�ccc�{{{�|||�rrr�rrr�rrr�yyy�~~~���������������������{{{�xxx�����aaaL      	   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ���Gvvv�"""�===�\\\�WWW�LLL�]]]�eee�nnn�ZZZ�^^^�fff������vvv�vvv�vvv�}}}�������������������������}}}���������bbbK         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ���Exxx�$$$�@@@�```�[[[�MMM�]]]�hhh�ppp�[[[�___�hhh���������yyy�zzz�zzz��������������������������������������fffF         ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��� ��� ���       ���Axxx�&&&�CCC�eee�___�MMM�```�jjj�sss�ZZZ�aaa�jjj���������}}}�~~~�~~~�����������������������������}}}���������uuu=         ��� ��� ��� ��� ��� ��� ���                   ��� ���    ���:����+++�FFF�jjj�bbb�MMM�aaa�jjj�sss�ZZZ�```�lll�������������������������������������������������{{{�������Ʀ���0   
   ��� ��� ��� ��� ��� ��� ��� ���             	         ���    ���#������������������������������������������������񴴴򓓓�zzz�yyy����������������������������������������gEEE      ��� ��� ��� ��� ��� ��� ��� ���    �|lp`T         	         %%%����¯Uհu~~}|�����������������xxx����J���:���3���0���1���2���2���4���<�����������������sssx���U���>���      ��� ��� ��� ��� ��� ��� ��� ��� ���    ��������LA9)         
         ϰ�D�L|�x gjif�������������nnn�MLG�   %                        eee�������������ggg�Y   *         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �����q��~���@700            Բ�S�Q�� z�x ujif�������������nnn�YSD� )            ���          eee�������������ggg�X   )         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� 湝F��A��n ��~��?5.2       ҭ�d�T��~ ��~ ��x �kif�������������nnn�eY@�S9 4C1      ��� ��� ���       fff�������������ggg�X   )         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� 깛N��6��l ��m ��~��<3,5ˣ�x�W��z ��{ ��| ��y �kif�������������nnn�n^>�wP @�e#��w   ��� ��� ���       ggg�������������ggg�X   )         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� 贕O��5��i ��l ��m ��~����Z��v ��x ��y ��z ��x �lie�������������nnn�xb;��bM��h9_[T	                  hhh�������������ggg�W   (         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� 豑O��3��f ��i ��k ��m ��u��r ��s ��u ��x ��x ��y�lie�������������nnn��g;���^iMH@   
               	   ggg�������������ggg�V   &         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� 欌P�2��d ��f ��i ��k ��m ��o ��r ��s ��u ��z��y�lid�������������uuu���f�3/)A   #                     !ccc�������������ggg�N   #      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� 橇P�~0��b ��d ��f ��i ��k ��m ��o ��r ��w��z	��y�}sh�����������������oon�M   :   1   -   ,   ,   -   0111Xjjj�������������ccc�   :         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� 䤂Q�z/��` ��b ��d ��f ��i ��k ��m ��t��x��x	��}ƚ~b꯯��������������www�nnn�\\\�[[[�[[[�[[[�[[[�[[[�aaa�bbb�����������������bbb�   0         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �~Q�x-��] ��` ��b ��d ��f ��i ��q
��t��u��w	���ц=ւ���������������������������|||�|||�|||�|||�{{{���������������������{{{�aaa�   #         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �yQ�v,��[ ��] ��` ��b ��d ��l��r��s��s��u
��~��+՜�������������������������������������������������������������������bbb�,         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �uQ�r*��Y ��[ ��] ��` ��j��o��o��q��q��r	��z����毟�r������������������������������������������������������������bbb�UUUo      
      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �rP�p)��V ��Y ��[ ��f��m��m��m��n��o��p	��v���0��֏��Y���ˀ���������������������������������������xxx�fff�bbb�CCC9      
      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �pK�o*��T ��V ��c��j��j��k��l��l��m��n	��q	��w���/��և�{MzzzG�uuu�lll�kkk�jjj�hhh�eee�ccc�eee�eee�LLL<               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ݍe!�~B��R ��`��g��h��h��i��j��k��k��l	��m��q��v���'�����}rl9RRR+++      
   
   
   
   
   
   	               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �`��b��e��e��f��g��g��h��i��i��j
��j��l��n��o�������ʁk\                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �h#�g��x;��g��d��d��f��f��f��h��h
��i��i��k��m��}����� e      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �}X	�en�g��i��l��o���q���t���w���y���|����������������綗.      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ������  ������  ���� ?  ����   ����   ����   ����   ����   ����   ����   ��     ��     ��     ��     ��     ��     ��    ��  �  ��  �  ��  �  ��  �  ��  �  ��  �  ��  �  ��  �  ��  �  ��  �  ��  �  ��  �  ����  ����  ����  ����  � ��  � ��  � ��  � ��  � ��  �   �  �   �  �   ��  � ��  � ��  � ���  � ���  � ?���  � ?���  � ���  (   @   �                              ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                       
                                                   	             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                               !   !                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                             "   $   &   (   )   +   ,   .   /   1   2   3   3   3   /   *   !            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           QqQ�ێS�蓇�葤�䎧�ጩ�ߋ������ߊ��݋��܊��ۉ��ډ��و��؈��ه�؆�~ԇ�n�u�AjF^   ;   1   #         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���        ��<����y�~�U�Y�E�H�E�H�E�H�E�H�E�H�E�H�E�H�E�I�E�I�E�I�E�I�E�I�E�I�E�I�H�M�h�o�����ڇ�+G   0         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���     �ի����e�h� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���n�t����:   '      
��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                �߫��N�Q� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���B�B�����s�z�   ,      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                              �ѡ��O�Q� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���>�>�C�C�h�k����   /      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                   �����O�Q� � � � � � � � � � � � � � � � � � � � � � � � � � ���:�:�?�?�B�B�P�P�����   /      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                    
                                                                     ZvZ�O�R� � � � � � � � � � � � � � � � � � � � � � ���6�6�;�;�?�?�B�B�F�F�����   /      ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                               :K:,���O�R� � � � � � � � � � � � � � � � � � ���2�2�7�7�;�;�>�>�B�B�F�F�����   .      ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                        )   .   1   2   2   2   2   2   2   2   2   2   2   2   2   2   2   2   2   2   2   2   2   3   3   57O7J���-�/� � � � � � � � � � � � � � ���/�/�3�3�7�7�;�;�>�>�B�B�F�F�����   ,      ��� ��� ��� ��� ��� ��� ��� ��� ��� ���          	   #3>F


I


J


J


J


J


J


J


J


J


J


J


J


J


J


J


J


J


J


J


J


J


J


K"R�̋�R�U��� � � � � � � � � � � � ���+�+�0�0�3�3�7�7�:�:�>�>�B�B�E�E�����   +      ��� ��� ��� ��� ��� ��� ��� ��� ���           """���F���o���������������������������������������������������������������������������������������������������������٬�S�V��� � � � � � � � � � � � ���'�'�,�,�/�/�3�3�7�7�:�:�>�>�B�B�E�E�����   *      ��� ��� ��� ��� ��� ��� ��� ��� ���           ���-���innn�^^^�\\\�ccc�iii�nnn�lll�hhh�aaa�WWW�ggg�sss����������������������������������������������������������X�Z����� � � � � � � � � � �
�
�#�#�(�(�,�,�/�/�3�3�6�6�:�:�>�>�A�A�E�E�����   )      ��� ��� ��� ��� ��� ��� ��� ��� ���           ���D����MMM��###�***�111�222�555�;;;�>>>�???�???�:::�999�888�888�===�===�>>>�<<<�===�@@@�BBB�EEE�GGG�NNN�s�t�L�M�����	�
��� � � � � � �	�	���$�$�(�(�+�+�/�/�3�3�6�6�:�:�>�>�A�A�E�E�����   '      ��� ��� ��� ��� ��� ��� ��� ��� ���           ���Fyyy�CCC��"""�)))�111�111�333�:::�>>>�>>>�>>>�:::�999�999�:::�AAA�BBB�BBB�@@@�AAA�DDD�FFF�III�NNN�k~l�L�M���������	�
��� � ����� � �$�$�(�(�+�+�/�/�2�2�6�6�:�:�=�=�A�A�E�E�����   &      ��� ��� ��� ��� ��� ��� ��� ��� ���           ���F}}}�FFF��"""�)))�111�000�222�:::�???�AAA�BBB�>>>�<<<�===�===�EEE�FFF�FFF�CCC�DDD�GGG�III�MMM�ana�J�K�)}*�%�&�!�"�������	�
������� � �#�#�'�'�+�+�/�/�2�2�6�6�:�:�=�=�A�A�D�D�����   %      ��� ��� ��� ��� ��� ��� ��� ��� ���           ���E����HHH��"""�)))�222�222�444�===�BBB�EEE�GGG�AAA�???�???�@@@�III�JJJ�KKK�HHH�HHH�JJJ�MMM�XaX�GxH�2t3�1|2�-�.�)�*�"�#������������� � �#�#�'�'�+�+�.�.�2�2�6�6�9�9�=�=�A�A�D�D�����   #      ��� ��� ��� ��� ��� ��� ��� ��� ���           ���E����JJJ��$$$�,,,�666�444�777�@@@�EEE�III�KKK�DDD�BBB�BBB�CCC�MMM�NNN�OOO�KKK�KKK�MMM�MRM�GiH�<l=�:s;�9{:�6�7�1�2�*�+�"�#� �!�$�%�#�$�$�%�"�#���#�#�'�'�,�,�.�.�2�2�6�6�9�9�=�=�@�@�D�D�����   !      
��� ��� ��� ��� ��� ��� ��� ��� ���           ���D����NNN��&&&�///�999�777�999�CCC�HHH�MMM�OOO�GGG�EEE�EEE�FFF�QQQ�SSS�SSS�OOO�OOO�PRP�J\J�FcG�DjE�CsD�AzB�?�@�:�;�2�3�-�.�0�1�+�,�(�)�,�-�+�,�#�$�#�#�)�)�߃�o�r�2�2�5�5�9�9�=�=�@�@�D�D�����         	��� ��� ��� ��� ��� ��� ��� ��� ���           ���D����MMM��'''�222�===�:::�<<<�EEE�KKK�PPP�SSS�JJJ�HHH�HHH�III�UUU�WWW�WWW�RRR�RRR�RSR�P[P�PdP�LiM�KqL�JzK�H�I�D�E�<�=�:�;�7�8�1�2�-�.�4�5�3�4�(�)�'�'�y�{�ꠡ���q�t�5�5�9�9�<�<�@�@�D�D�����         ��� ��� ��� ��� ��� ��� ��� ��� ���           ���C����HHH��)))�444�@@@�<<<�===�HHH�MMM�SSS�WWW�MMM�JJJ�KKK�KKK�YYY�ZZZ�[[[�VVV�WWW�VVV�XYX�XcX�ThT�TqU�U{V�S�T�P�Q�H�I�A�B�?�@�8�9�4�5�<�=�<�=�0�0�s�u�ޜ�+v�v����t�v�8�8�<�<�@�@�D�D�����         ��� ��� ��� ��� ��� ��� ��� ��� ���           ���Czzz�DDD��+++�777�DDD�???�???�JJJ�PPP�UUU�[[[�QQQ�MMM�MMM�MMM�]]]�___�___�YYY�YYY�YYY�[[[�`a`�\g\�]q]�_|`�^�_�[�\�Q�R�K�L�G�H�?�@�;�<�E�F�G�H�w�y�ʔ�      �ɏ����v�x�<�<�@�@�F�G�����      
   ��� ��� ��� ��� ��� ��� ��� ��� ���           ���Bqqq�@@@��---�:::�GGG�AAA�@@@�LLL�RRR�XXX�^^^�SSS�OOO�OOO�PPP�aaa�bbb�ccc�]]]�^^^�]]]�^^^�ddd�fgf�grg�j~j�i�j�g�h�Z�[�T�U�P�Q�F�G�B�C�N�O��ȃ��ͫ�-      	      ������x�z�@�@�Z�[�����         ��� ��� ��� ��� ��� ��� ��� ��� ���           ���Bmmm�@@@��...�===�KKK�DDD�BBB�NNN�SSS�ZZZ�aaa�VVV�RRR�QQQ�SSS�eee�fff�ggg�```�```�```�aaa�ggg�iii�pqp�v�v�v�v�s�t�f�g�]�^�X�Y�N�O�J�K�z�|��κ圞�x   *      	         ������{�~��������         ��� ��� ��� ��� ��� ��� ��� ��� ���           ���Avvv�DDD��111�???�OOO�FFF�CCC�OOO�VVV�\\\�bbb�XXX�TTT�SSS�TTT�hhh�jjj�kkk�ccc�ccc�ddd�ddd�jjj�mmm�ttt�������������s�t�g�h�b�c�W�X�k�l��������ۜ��w   *      	             �����Ȥ���ێ         ��� ��� ��� ��� ��� ��� ��� ��� ���           ���A}}}�III�   �111�BBB�SSS�HHH�EEE�RRR�XXX�^^^�eee�[[[�UUU�UUU�VVV�kkk�nnn�nnn�fff�ggg�ggg�fff�mmm�ppp�xxx���������������r�s�m�n�m�n����������ޛ��w   *      	      ���         �����:              ��� ��� ��� ��� ��� ��� ��� ��� ���           ���@����OOO�!!!�444�EEE�VVV�III�EEE�TTT�ZZZ�```�hhh�]]]�WWW�XXX�XXX�ppp�qqq�rrr�iii�jjj�kkk�jjj�ppp�sss�{{{�����������������|�|�|�|���vvv�|||����ᛛ�w   *      	      ��� ��� ���                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           ���@����PPP�!!!�555�HHH�ZZZ�LLL�FFF�TTT�[[[�bbb�jjj�^^^�YYY�YYY�[[[�rrr�uuu�vvv�mmm�mmm�mmm�lll�sss�uuu��������������������������|||�www�ttt����䚚�v   *      	      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           ���@����QQQ�###�777�JJJ�___�NNN�GGG�VVV�]]]�ddd�jjj�^^^�[[[�ZZZ�\\\�vvv�yyy�yyy�ooo�ppp�ppp�ppp�vvv�xxx������������������������������xxx�nnn����皚�v   *      	      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           ���@����QQQ�"""�999�MMM�ccc�PPP�HHH�YYY�___�fff�mmm�___�]]]�]]]�]]]�yyy�|||�}}}�rrr�sss�sss�sss�yyy�zzz���������������������������������{{{�xxx����晙�t   )      	      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           ���@����RRR�###�;;;�PPP�ggg�RRR�HHH�YYY�```�ggg�ooo�___�]]]�]]]�___�|||���������vvv�vvv�vvv�uuu�|||�|||���������������������������������|||��������⚚�t   (            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           ���=����SSS�$$$�===�RRR�kkk�TTT�III�[[[�aaa�iii�ppp�```�]]]�___�___�������������xxx�yyy�yyy�yyy�����������������������������������������~~~��������ݛ��q   &            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           ���;����SSS�%%%�???�UUU�ppp�VVV�III�[[[�ccc�jjj�qqq�```�^^^�aaa�bbb�������������zzz�{{{�{{{�{{{�������������������������������������������������آ��l   "             ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                      ��� ���           ���8����TTT�'''�AAA�XXX�ttt�YYY�III�\\\�ccc�jjj�sss�```�\\\�aaa�ccc�������������}}}�~~~�������������������������������������������|||��������ѭ��d                ��� ��� ��� ��� ��� ��� ��� ��� ���                                        ���6����^^^�(((�DDD�[[[�yyy�ZZZ�III�]]]�eee�lll�sss�aaa�\\\�```�ccc������������������������������������������������������������������zzz�������ü���[      	      ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                      ���%���Y����aaa�nnn�������������qqq�������������������������������������������������yyy�nnn�zzz����������������������������������������������������z���?             ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                   
                  ������@���\�������ݠ��𞞞������������������������㵵�к����������������������ů��Π��ԑ��ܒ��ۢ��թ��𳳳������������������������ݼ����������y���^{{{             ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ɫ�7            	                  	���"�ūd׫f}��l�xxx�����������������rrr�mmm�___F~~~7���+���&���$���#���#���#���$���$���&���+~~~�������������������ppp�ccc~dddR���?���*   
             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��}�˦�����
            	            	&"���a�J~�z f�rU�kkk�����������������bbb�RPM�   /                                 ggg�ttt�����������������\\\�000j   6   !                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �Þ���4���_�给�	%               
   )%!�ßp�N�ـ s�z p�sS�kkk�����������������bbb�ZUK� 3                                   	hhh�vvv�����������������\\\�000j   6                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �Ǣ��o��p ���_�乗�
	(             �Þ��O�� ��~ ~�y z�tQ�kkk�����������������bbb�`YH�<* ;'                  ��� ���          	hhh�www�����������������\\\�000j   5                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �xe�����l ��n ��p ���_�㸗�
	)   "   �����P��~ ��~ ��} ��y ��tP�kkk�����������������bbb�h]F�W; DV< )D0             ��� ���          	hhh�yyy�����������������\\\�000j   5                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��s�����k ��l ��n ��o ���`�ⷖ�
,*罚��Q��z ��{ ��| ��| ��y ��tN�kkk�����������������bbb�n`E�oK LwQ 1�^	��x          ��� ���          	hhh�{{{�����������������\\\�000j   5                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��l�����h ��j ��k ��m ��o ���`�ⷖ�滙��S��w ��y ��y ��z ��z ��y ��uM�kkk�����������������bbb�tbC��U S�a:��Z4���                           	ggg�}}}�����������������\\\�000i   5                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��j�����f ��h ��j ��k ��m ��o ���`���T��t ��u ��w ��x ��x ��y ��x ��uL�kkk�����������������bbb�ydA��\ \��TW���-                        ggg�{{{�����������������\\\�111h   4                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �g�����e ��f ��h ��j ��k ��m ��o ��q ��s ��s ��u ��w ��x ��x ��z��vK�kkk�����������������bbb�~f?���P|��vJ                        
   fff�ttt�����������������\\\�111h   2                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �}e�����c ��e ��f ��h ��j ��k ��m ��o ��q ��r ��s ��u ��v ��{��z��uI�kkk�����������������eee��a}ik   ,                              eee�nnn�����������������\\\�222e   /                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �w_��~��a ��c ��e ��f ��h ��j ��k ��m ��o ��q ��r ��s ��y��{��z��w3�fff�����������������sss�yvr�K   :   .   '   #   "   !   !   "   #   &   -ccc�sss�����������������]]]�E   +      
      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �u]��{��` ��a ��c ��e ��f ��h ��j ��k ��m ��o ��q ��v��y
��z��{
���jii���������������������nnn�***`N   B   <   9   8   8   8   8   9   <K___���������������������aaa�   :   %             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �s[��x��^ ��` ��a ��c ��e ��f ��h ��j ��k ��m ��t	��x��x
��x	��}���usq���������������������www�lll�kkk�```�___�```�```�```�```�```�```�bbb�^^^�nnn�����������������zzz�bbb�   2                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �nV��u��\ ��^ ��` ��a ��c ��e ��f ��h ��j ��q
��u��v��w
��x��~��ʉ}q�����������������������������}}}�rrr�nnn�nnn�nnn�nnn�nnn�nnn�nnn�uuu�������������������������ccc�^^^�   (      
      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �lS��r��Z ��\ ��^ ��` ��a ��c ��e ��f ��n��s��s��t��u
��x��~�����6�~}|�������������������������������������������������������������������������������������xxx�aaa�   -               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �jQ��o��Y ��Z ��\ ��^ ��` ��a ��c ��l��p��q��r��r��s
��v��}�� ����Ღ�ؕ�����������������������������������������������������������������������������������^^^�HHHc         	          ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �iO��l��W ��Y ��Z ��\ ��^ ��` ��i��n��o��o��p��q��q
��t��z���N��ϳ�~~}T���ۘ�����������������������������������������������������������������������vvv�^^^�bbb�         
          ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �oS�i��U ��W ��Y ��Z ��\ ��g��m��m��m��n��n��o��p
��q
��w��}���w��Ī��T����������������������������������������������������������������yyy�ccc�bbb�MMMV         
             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �rT�g��S ��U ��W ��Y ��d��j��k��l��l��l��m��m��n
��o	��r��x��~���w��ũ�xwwL���M����{{{�rrr�ggg�^^^�\\\�\\\�\\\�\\\�\\\�\\\�\\\�^^^�bbb�eee�eee�                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� uL7��j��R ��S ��U ��b��i��i��i��j��k��k��l��l��l��m	��n��r��x��|���s��ŧ�mkj?jjj5lll-ddd$HHH""""""""""""                                        ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��jݿT��R ��`��g��g��h��h��h��i��j��j��k��l��k	��l��n��q
��v��y���m��ä�[ZX,RRR>>>      	                                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �f~�{>��^��e��e��f��f��g��g��h��h��i��i��j��k	��k��k��n��o��q��u���h��ģ�0,*                                                    ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    f@-��l��~E��d��d��d��e��e��f��f��g��g��h��h��i
��j��j��k��m��m��o ��q ���y��Ȧ�                                                       ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���        у]��j��k���P��|=��|<��|;��}:��~:��9��8��8��8��7��7���6���6���5���5���K���z��Ü�ߵ�)             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           �f#��pZ��m��o��q��t���v���y���{���~��������������������������������j칙5                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �����������������������������  �����  �����  �����  �����  �����  ������ ������ ������ ������ ��     ��     ��     ��     ��     ��     ��     ��     ��     ��    ��    ��    ?��    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ����   ��������������������������� ����� ����  ����  ����  ����  ����  ����  ����    ���    ���    ���    ?���   ?���   ����  ���� ������ ������  ������  �����  ������ �����(   �                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                	   	   	   
   
   
   
                                                                        
   	                            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                    	                                                                                                               	                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                 
                                                                                                                           	                   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                  !   !   "   "   #   #   $   $   %   %   %   %   $   #   "                         	               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                              
                               !   "   #   #   $   %   %   &   &   '   (   (   )   *   *   +   ,   ,   -   .   .   /   /   /   .   -   ,   *   '   #                  
            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                               	                         "   $   %   '   (   )   *   +   ,   ,   -   .   /   /   0   1   2   3   3   4   5   6   6   7   8   8   8   8   7   6   3   0   ,   (   "               	         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                              
         1S7%X�\:T�X=P�T?M{QBKxODIuMFHtLFGrKGFpIIEnHJDmHKDmHKClGLCkFMBiEMAhDN@gDO@fCP?eBQ>dAR>cAS>cAS<a?T<`?U<`?U;_>V;^=W:]=X:]=X0J   @   ?   >   <   9   5   0   *   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                           ~Ƅ+��x�������ܝ������������������������������������������������������������������������������������������������������������������������������ݒ�u�|�CnHd   A   =   8   1   +   #            
      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                      @`@���m��������������������������������������������������������������������������������������������������������������������������������������������������������}ʄ�H   ?   8   1   )   !            	   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���               ��+�����������^�b�3�5��� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���7�;�_�f������������JwOg   >   7   /   &            
   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���        �������������#�%� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �"�$�������������BjE`   ;   3   *   !            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���            ���<���Ǔ��M�O� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��������������A   7   .   $            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���           ���=���Ȕ��L�O� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �
�
�<�<�I�I���������yƃ�   :   0   '            	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���               ���=���Ȕ��L�O� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �
�
�:�:�B�B�D�D�b�d���������6Y9Q   2   (            
��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                                                                                                    ���=���ɔ��L�O� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �	�	�8�8�@�@�B�B�D�D�F�F���������l�t�   3   *             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                                                                             ��@���ɔ��M�O� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �	�	�6�6�>�>�@�@�B�B�D�D�E�E�z�}������Ս�   4   *   !         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                                                                                     ��A���˔��M�O� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �	�	�5�5�<�<�>�>�@�@�B�B�C�C�E�E�b�d��������   4   +   !         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                                                                                              ��C���˔��M�O� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���3�3�:�:�<�<�>�>�@�@�B�B�C�C�E�E�L�L���������   4   +   !         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                      	   	   	   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
         �؛G���͔��M�O� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���1�1�8�8�:�:�<�<�>�>�@�@�A�A�C�C�E�E�G�G���������   4   *   !         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                             	                                                                                                                                                         �˒K���ϔ��M�P� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���0�0�6�6�8�8�:�:�<�<�>�>�@�@�A�A�C�C�E�E�G�G���������   3   *   !         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                           	                                                                                                                                                                  ���Q���є��M�P� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���.�.�4�4�6�6�8�8�:�:�<�<�>�>�?�?�A�A�C�C�E�E�G�G���������   3   *   !         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                       	                               !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   !   "   #   #   %v�|[���ӓ��M�P� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���,�,�2�2�4�4�6�6�8�8�:�:�<�<�>�>�?�?�A�A�C�C�E�E�G�G���������   2   )             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                        	                  #   &   (   *   +   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   ,   -   -   .   /   1k�pd��ה��M�P� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ���*�*�1�1�2�2�4�4�6�6�8�8�:�:�<�<�=�=�?�?�A�A�C�C�E�E�F�F���������   1   (             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                    	               #   (   -   0   3   5   6   7   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   8   9   9   :   ;FdIW��˔��b�e��� � � � � � � � � � � � � � � � � � � � � � � � � � � � ���)�)�/�/�1�1�2�2�4�4�6�6�8�8�:�:�<�<�=�=�?�?�A�A�C�C�E�E�F�F���������   1   (            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                $   +   1   7   ;   >   @   A   B   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   C   D   D   D   D   E?XB]�ߥÐ��]�`��� � � � � � � � � � � � � � � � � � � � � � � � � � � � ���'�'�-�-�/�/�0�0�2�2�4�4�6�6�8�8�:�:�;�;�=�=�?�?�A�A�C�C�D�D�F�F���������   0   '            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	         "&&&1###9!!!@FJNPRSSSSSSSSSSSSSSSSSSSTTTTTTTTTTTTTTTTTTTTTTTTUUUL]Li�ڥ����Y�[��� � � � � � � � � � � � � � � � � � � � � � � � � � � � ���%�%�+�+�-�-�/�/�0�0�2�2�4�4�6�6�8�8�:�:�;�;�=�=�?�?�A�A�C�C�D�D�F�F���������   /   '            
��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                    
   WWW ���Q���k���v���|������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������אߔ�V�X��� � � � � � � � � � � � � � � � � � � � � � � � � � � � ���#�#�)�)�+�+�-�-�.�.�0�0�2�2�4�4�6�6�8�8�9�9�;�;�=�=�?�?�A�A�B�B�D�D�F�F���������   .   &            
��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                    ��� ���a���k���r���|�������ڊ��݌��ގ��ݒ��ޔ��ݗ��ܙ��ܖ��ۖ��ܕ��ݔ��ޓ��ߑ������⍍�㑑�����ߘ��ݛ��ܞ��ڡ��ئ��֧��ԧ��է��է��ԩ��ԩ��Ԫ��ө��ө��ԩ��ԩ��ԩ��ԩ��ԩ��Ԫ��ԫ��ԫ��ԫ��Ԭ��ԭ��ԭ��Ԯ��ӯ��ӯ��ӱ��Բ��Գ��Է��ڿ���ܕ�X�Z�	�
��� � � � � � � � � � � � � � � � � � � � � � � � � � ���!�!�'�'�)�)�+�+�-�-�.�.�0�0�2�2�4�4�6�6�8�8�9�9�;�;�=�=�?�?�A�A�B�B�D�D�F�F���������   -   %            
��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 ���S���f���m����hhh�ccc�fff�jjj�mmm�qqq�uuu�yyy�|||������}}}�zzz�www�sss�lll�fff�^^^�ccc�mmm�vvv���������������������������������������������������������������������������������������������������������������������������׿��֓�Z�\��������� � � � � � � � � � � � � � � � � � � � � � ��� � �%�%�'�'�)�)�+�+�,�,�.�.�0�0�2�2�4�4�6�6�7�7�9�9�;�;�=�=�?�?�@�@�B�B�D�D�F�F���������   -   %            
��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 ������a���f����\\\�[[[�]]]�LLL�KKK�NNN�PPP�TTT�WWW�YYY�\\\�\\\�\\\�[[[�\\\�[[[�ZZZ�YYY�UUU�UUU�YYY�___�bbb�ccc�fff�iii�lll�nnn�nnn�nnn�rrr�rrr�rrr�rrr�rrr�qqq�ppp�qqq�qqq�rrr�sss�ttt�uuu�uuu�www�xxx�yyy�zzz�|||�}}}�~~~����������Ƈ�V�W�������	�
����� � � � � � � � � � � � � � � � � � �����#�#�%�%�'�'�)�)�+�+�,�,�.�.�0�0�2�2�4�4�6�6�7�7�9�9�;�;�=�=�>�>�@�@�B�B�D�D�F�F���������   ,   $            
��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���+���a���gmmm�UUU�JJJ���!!!�%%%�'''�,,,�000�222�333�000�333�666�:::�===�???�>>>�???�>>>�???�???�<<<�999�999�999�888�888�888�888�<<<�===�===�===�===�<<<�:::�;;;�<<<�===�???�@@@�@@@�AAA�DDD�EEE�EEE�GGG�JJJ�KKK�WZW�����u�v�P�R����������	������� � � � � � � � � � � � � � �����!�!�#�#�%�%�'�'�)�)�*�*�,�,�.�.�0�0�2�2�4�4�5�5�7�7�9�9�;�;�=�=�>�>�@�@�B�B�D�D�F�F���������   +   #            	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���.���a���gddd�[[[�(((���!!!�%%%�'''�,,,�///�111�333�000�222�666�:::�<<<�>>>�>>>�>>>�>>>�???�???�<<<�999�999�888�888�777�777�777�===�>>>�>>>�???�???�???�===�===�>>>�???�@@@�AAA�CCC�CCC�EEE�GGG�HHH�III�LLL�VXV����q�s�N�P�������������	�
������� � � � � � � � � � �������!�!�#�#�%�%�'�'�)�)�*�*�,�,�.�.�0�0�2�2�4�4�5�5�7�7�9�9�;�;�<�<�>�>�@�@�B�B�D�D�F�F���������   *   #            	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���-���a���gddd�___����   �$$$�'''�,,,�///�111�222�///�222�555�999�;;;�===�>>>�>>>�???�>>>�>>>�;;;�888�888�999�888�888�999�999�???�@@@�AAA�AAA�AAA�AAA�???�???�@@@�AAA�BBB�CCC�EEE�EEE�HHH�HHH�JJJ�LLL�VWV�z�z�m�n�N�O�����������������	�
������� � � � � � ���������!�!�#�#�%�%�'�'�(�(�*�*�,�,�.�.�0�0�2�2�3�3�5�5�7�7�9�9�;�;�<�<�>�>�@�@�B�B�D�D�F�F���������   *   #            	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���.���`���ghhh�bbb����   �$$$�&&&�,,,�///�111�222�///�111�555�999�;;;�===�>>>�>>>�>>>�>>>�???�<<<�999�999�:::�:::�:::�:::�;;;�AAA�BBB�CCC�DDD�CCC�CCC�@@@�AAA�AAA�CCC�DDD�EEE�FFF�GGG�III�KKK�LLL�TUT�t}u�g�h�L�M�$�%� �!�� ���������������	�
������� � �����������!�!�#�#�%�%�'�'�(�(�*�*�,�,�.�.�0�0�2�2�3�3�5�5�7�7�9�9�:�:�<�<�>�>�@�@�B�B�D�D�F�F���������   )   "            	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���.���`���glll�fff����   �$$$�&&&�,,,�///�111�222�...�111�444�888�:::�===�???�???�@@@�AAA�AAA�>>>�;;;�;;;�;;;�;;;�<<<�<<<�<<<�CCC�DDD�EEE�EEE�EEE�EEE�BBB�BBB�CCC�DDD�EEE�GGG�HHH�III�KKK�MMM�RSR�nsn�b�c�J�K�(|)�&~'�$�%�#�$�!�"���������������	�
�����������������!�!�#�#�%�%�&�&�(�(�*�*�,�,�.�.�0�0�1�1�3�3�5�5�7�7�9�9�:�:�<�<�>�>�@�@�B�B�D�D�E�E���������   (   !            	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���.���`���gppp�hhh����   �$$$�&&&�,,,�///�111�222�...�000�555�888�<<<�>>>�AAA�BBB�BBB�CCC�DDD�@@@�===�>>>�===�===�===�>>>�>>>�EEE�FFF�GGG�GGG�GGG�GGG�EEE�EEE�EEE�EEE�GGG�HHH�III�KKK�MMM�RSR�hkh�\�]�I�J�-x.�+{,�*~+�'(�'�(�$�%�"�#���������������	�
�	�
�������������!�!�#�#�%�%�&�&�(�(�*�*�,�,�.�.�0�0�1�1�3�3�5�5�7�7�8�8�:�:�<�<�>�>�@�@�B�B�D�D�E�E���������   (   !            	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���.���`���fuuu�mmm�����###�&&&�---�000�222�333�///�222�555�:::�===�???�BBB�DDD�EEE�FFF�FFF�BBB�>>>�???�???�???�>>>�???�???�GGG�HHH�III�III�JJJ�III�GGG�GGG�GGG�GGG�III�III�KKK�LLL�RRR�bdb�WzX�H�I�3t4�0w1�/z0�/0�+,�+�,�(�)�&�'�"�#�����������������������������!�!�#�#�$�$�&�&�(�(�*�*�,�,�.�.�/�/�1�1�3�3�5�5�7�7�8�8�:�:�<�<�>�>�@�@�B�B�C�C�E�E���������   '                	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���.���_���fxxx�ppp����   �$$$�&&&�...�222�444�555�000�333�888�<<<�???�AAA�DDD�EEE�GGG�GGG�GGG�DDD�@@@�@@@�@@@�@@@�@@@�AAA�AAA�III�KKK�KKK�KKK�LLL�KKK�III�HHH�JJJ�III�JJJ�LLL�MMM�NNN�Z[Z�RqS�FxG�6o7�5s6�3u4�3z4�2}3�/0�/�0�,�-�*�+�&�'�!�"�������������������� �������!�!�"�"�$�$�&�&�(�(�*�*�,�,�.�.�/�/�1�1�3�3�5�5�6�6�8�8�:�:�<�<�>�>�@�@�B�B�C�C�E�E���������   &               	��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���.���_���f}}}�ttt����   �%%%�(((�///�333�666�777�111�444�888�===�@@@�CCC�EEE�HHH�HHH�III�JJJ�EEE�AAA�BBB�BBB�AAA�BBB�BBB�CCC�LLL�MMM�MMM�NNN�MMM�NNN�JJJ�JJJ�JJJ�JJJ�KKK�MMM�NNN�STS�LeM�DnE�;k<�9n:�9r:�7u8�7y8�7~8�3~4�3�4�1�2�.�/�*�+�%�&�"�#�� �����#�$�"�#�!�"� �!�� �#�$�"�#�����!�!�"�"�$�$�&�&�(�(�*�*�,�,�-�-�/�/�1�1�3�3�5�5�6�6�8�8�:�:�<�<�>�>�@�@�A�A�C�C�E�E���������   %               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���-���_���e����xxx����!!!�&&&�)))�111�555�777�888�222�666�:::�???�AAA�DDD�GGG�JJJ�KKK�KKK�KKK�GGG�CCC�CCC�CCC�CCC�DDD�DDD�EEE�MMM�OOO�OOO�OOO�OOO�OOO�LLL�MMM�LLL�LLL�MMM�NNN�PPP�G[G�DfE�@fA�>i?�=m>�=r>�;t<�;y<�;}<�89�8�9�5�6�2�3�.�/�)�*�&�'�#�$�!�"�(�)�'�(�%�&�$�%�#�$�!�"�)�*�&�'�"�#� �!� � �"�"�$�$�&�&�(�(�*�*�3�3�-�-�/�/�1�1�3�3�4�4�6�6�8�8�:�:�<�<�>�>�@�@�A�A�C�C�E�E���������   $               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���-���^���e����{{{����"""�'''�***�222�777�999�:::�333�777�:::�@@@�CCC�FFF�HHH�KKK�MMM�MMM�NNN�JJJ�DDD�EEE�EEE�DDD�EEE�EEE�EEE�OOO�QQQ�QQQ�RRR�RRR�RRR�NNN�NNN�NNN�NNN�NNN�PPP�JXJ�E^E�FcG�DfE�CiD�AlB�AqB�?t@�@yA�?}@�<~=�=�>�9�:�6�7�2�3�,�-�*�+�'�(�-�.�,�-�*�+�(�)�'�(�%�&�$�%�.�/�+�,�%�&�$�%�!�"�"�"�$�$�&�&�(�(�5�5����n�q�/�/�1�1�3�3�4�4�6�6�8�8�:�:�<�<�>�>�?�?�A�A�C�C�E�E���������   #               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���-���^���d����|||����###�(((�+++�444�999�;;;�<<<�444�777�<<<�AAA�DDD�GGG�JJJ�MMM�NNN�OOO�PPP�KKK�FFF�FFF�EEE�EEE�FFF�FFF�GGG�QQQ�SSS�TTT�TTT�TTT�TTT�PPP�PPP�PPP�PPP�PPP�MTM�JZJ�I]I�IbI�IfJ�FhG�FlG�FqG�CsD�CxD�D}E�@~A�A�B�>�?�<�=�7�8�0�1�/�0�2�3�1�2�0�1�-�.�+�,�)�*�(�)�'�(�3�4�0�1�(�)�&�'�"�#�"�#�$�$�&�&�2�3�����������o�r�1�1�2�2�4�4�6�6�8�8�:�:�<�<�>�>�?�?�A�A�C�C�E�E���������   !               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���-���^���d����|||����$$$�)))�,,,�666�:::�<<<�===�555�888�<<<�BBB�FFF�III�LLL�NNN�QQQ�QQQ�RRR�MMM�GGG�GGG�GGG�GGG�GGG�GGG�HHH�SSS�UUU�VVV�VVV�VVV�VVV�RRR�RRR�QQQ�RRR�RSR�PVP�NYN�N^N�NbN�MfM�JgK�IkJ�JpK�HsI�GwH�H}I�E~F�G�H�C�D�@�A�<�=�6�7�8�9�7�8�5�6�4�5�1�2�.�/�,�-�+�,�*�+�7�8�6�7�+�,�)�*�$�%�#�$�$�%�1�1�������������ئ���q�s�2�2�4�4�6�6�8�8�:�:�<�<�=�=�?�?�A�A�C�C�E�E���������               
   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���-���]���d����xxx����$$$�+++�---�777�<<<�>>>�???�666�999�>>>�CCC�GGG�III�LLL�OOO�RRR�SSS�SSS�NNN�HHH�III�HHH�III�III�III�III�VVV�WWW�WWW�YYY�XXX�WWW�SSS�SSS�TTT�TTT�TTT�STS�SYS�Q\Q�RbR�PdP�NgN�MjN�NpO�MsN�MxN�M}N�I~J�L�M�H�I�E�F�A�B�>�?�=�>�;�<�9�:�8�9�5�6�1�2�/�0�.�/�-�.�=�>�:�;�.�/�,�-�&�'�$�%�/�0��ۇ�����KpK�ݜJ���ا���r�t�4�4�6�6�8�8�:�:�;�;�=�=�?�?�A�A�C�C�D�D���������               
   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���-���]���dyyy�rrr����%%%�,,,�...�999�>>>�@@@�AAA�666�:::�???�EEE�HHH�KKK�NNN�QQQ�SSS�VVV�VVV�PPP�JJJ�JJJ�JJJ�JJJ�KKK�KKK�KKK�WWW�YYY�ZZZ�YYY�ZZZ�ZZZ�UUU�UUU�UUU�UUU�VVV�UUU�VWV�V\V�VaV�VfV�SgS�QjQ�SpT�QsR�RxS�S~T�N~O�Q�R�N�O�J�K�H�I�B�C�@�A�?�@�=�>�<�=�8�9�5�6�3�4�1�2�0�1�A�B�?�@�1�2�0�1�'�)�.�/�؄���ګ�HcH      
��F���ק���s�u�6�6�8�8�:�:�;�;�=�=�?�?�A�A�C�C�D�D���������               	   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���-���]���dsss�mmm����&&&�---�000�;;;�@@@�BBB�BBB�777�:::�???�FFF�JJJ�LLL�OOO�RRR�VVV�WWW�XXX�RRR�LLL�LLL�KKK�KKK�LLL�LLL�LLL�YYY�[[[�[[[�\\\�\\\�[[[�VVV�VVV�WWW�VVV�XXX�WWW�XXX�XYX�Z`Z�YdY�VfV�WkW�XqX�UrV�VxW�X~Y�TU�W�X�T�U�R�S�N�O�F�G�D�E�C�D�A�B�@�A�;�<�8�9�6�7�5�6�3�4�F�G�C�D�5�6�3�4�3�4�ԁ���ԫ宔@O@             ��D���ب���t�w�8�8�9�9�;�;�=�=�?�?�A�A�B�B�D�D���������                  ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���,���\���cmmm�ggg����&&&�...�111�<<<�BBB�DDD�DDD�888�<<<�AAA�FFF�KKK�NNN�PPP�SSS�WWW�ZZZ�ZZZ�TTT�LLL�MMM�LLL�LLL�MMM�MMM�NNN�[[[�]]]�]]]�^^^�^^^�^^^�YYY�XXX�YYY�YYY�YYY�XXX�ZZZ�[[[�^_^�]c]�[f[�ZjZ�[o[�ZsZ�[x\�]^�YZ�\�]�Z�[�W�X�S�T�K�L�I�J�G�H�F�G�D�E�?�@�;�<�:�;�8�9�7�8�K�L�I�J�8�9�@�A�|�~�ܝΧڪ�.B.'         	         ���D���٩���v�x�9�9�;�;�=�=�?�?�A�A�B�B�D�D���������            	      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���,���\���cfff�aaa����'''�///�222�===�DDD�EEE�EEE�999�===�AAA�HHH�LLL�OOO�QQQ�TTT�WWW�[[[�]]]�UUU�MMM�NNN�NNN�NNN�NNN�OOO�OOO�\\\�___�___�```�___�```�ZZZ�ZZZ�ZZZ�ZZZ�ZZZ�ZZZ�[[[�]]]�aaa�aba�`f`�_j_�aqa�^r^�`y`�d�e�_�`�b�c�`�a�]�^�W�X�O�P�M�N�L�M�J�K�G�H�B�C�?�@�=�>�<�=�:�;�R�S�M�N�D�E�Ѐ�۟Рͤ�&1&/                        ���C���٩���w�z�;�;�=�=�?�?�@�@�B�B�N�N���������                  ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���,���\���b___�[[[����(((�000�222�???�EEE�GGG�HHH�999�>>>�BBB�JJJ�LLL�PPP�SSS�VVV�YYY�\\\�^^^�VVV�NNN�OOO�OOO�OOO�OOO�OOO�PPP�^^^�aaa�```�bbb�aaa�aaa�\\\�\\\�\\\�]]]�]]]�\\\�\\\�^^^�ccc�eee�efe�bhb�fqf�csc�eye�i�i�d�e�h�i�f�g�c�d�]�^�S�T�R�S�P�Q�N�O�L�M�F�G�B�C�A�B�?�@�>�?�U�V�X�Y�~΀�ݩܬί�% 7   %                           ���C���٪���x�z�=�=�?�?�@�@�B�B�d�f���������         	         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���,���\���bXXX�UUU���   �)))�111�444�AAA�GGG�III�III�:::�>>>�CCC�KKK�NNN�QQQ�TTT�VVV�ZZZ�]]]�___�XXX�PPP�QQQ�PPP�OOO�PPP�PPP�PPP�```�bbb�ccc�ddd�ddd�ddd�^^^�^^^�^^^�^^^�^^^�___�^^^�```�ddd�fff�fff�ghg�jpj�iti�jzj�n�n�j�j�o�p�m�n�i�j�c�d�Y�Z�W�X�U�V�R�S�P�Q�J�K�F�G�D�E�C�D�A�B�`�a��ˆ��ק���Ży{y`   0   %                              ���C���ګ���z�|�>�>�@�@�B�B�|�~���������   
   	            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���,���[���bRRR�SSS���   �)))�111�444�BBB�III�KKK�JJJ�:::�???�DDD�KKK�OOO�RRR�UUU�XXX�[[[�___�aaa�ZZZ�QQQ�RRR�PPP�QQQ�PPP�RRR�RRR�bbb�ddd�fff�fff�fff�eee�___�___�___�___�```�___�```�aaa�eee�hhh�hhh�jjj�opo�ntn�p{p�t�t�o�o�t�t�s�t�n�o�j�k�_�`�\�]�Z�[�W�X�U�V�O�P�I�J�H�I�F�G�H�I��ǈ��Ӯ���º����qqq[   0   %                                  ���C���۫���{�}�@�@�D�D����������U                  ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���,���[���aYYY�XXX���   �***�333�555�DDD�KKK�MMM�MMM�;;;�???�DDD�LLL�PPP�SSS�VVV�YYY�\\\�___�ccc�[[[�QQQ�RRR�RRR�RRR�RRR�SSS�SSS�ddd�fff�ggg�ggg�hhh�ggg�aaa�aaa�aaa�aaa�aaa�aaa�aaa�bbb�fff�iii�iii�lll�qqq�sts�tzt�z�z�u�u�|�|�y�y�v�w�o�p�d�e�a�b�^�_�[�\�Z�[�S�T�M�N�L�M�M�N�p�q��ɨ�������������rrrZ   /   $                                      ���B���ڬ���|�~�t�v���������g�g                  ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���,���[���a___�^^^���   �+++�444�777�FFF�MMM�OOO�NNN�;;;�@@@�EEE�MMM�QQQ�TTT�XXX�ZZZ�]]]�aaa�ddd�]]]�SSS�SSS�SSS�SSS�TTT�TTT�UUU�eee�iii�jjj�iii�jjj�iii�bbb�ccc�ccc�bbb�ccc�ccc�ccc�ccc�hhh�jjj�lll�nnn�sss�uuu�{|{�����|�|�������{�{�v�w�i�j�f�g�c�d�`�a�_�`�W�X�Q�R�Q�R�m�n���������������������qqqY   /   $                     ��� ���              ���B���ۭ�������������D                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���+���Z���afff�ddd���   �+++�444�888�GGG�NNN�QQQ�PPP�<<<�@@@�GGG�NNN�RRR�UUU�YYY�[[[�^^^�bbb�eee�^^^�TTT�UUU�TTT�TTT�UUU�UUU�UUU�ggg�kkk�jjj�kkk�kkk�kkk�ddd�ddd�eee�eee�eee�ddd�fff�eee�jjj�lll�mmm�ooo�ttt�vvv����������������������}�}�n�o�k�l�i�j�e�f�d�e�Z�[�W�X�l�m�������������������������qqqY   /   $                     ��� ���                  ���B���ۨ������                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���+���Z���ammm�jjj���!!!�,,,�666�999�HHH�QQQ�QQQ�QQQ�===�@@@�GGG�OOO�RRR�VVV�YYY�]]]�```�ccc�ggg�___�UUU�UUU�VVV�TTT�UUU�UUU�VVV�iii�lll�mmm�mmm�mmm�lll�fff�eee�fff�fff�eee�fff�fff�fff�kkk�mmm�nnn�qqq�vvv�xxx�����������������������������t�t�p�q�m�n�k�l�i�j�a�b�l�m�}�~�����rsr�����������������qqqY   /   $                     ��� ��� ���                   ���B���Ġ�                           ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���+���Z���asss�ppp���!!!�---�777�:::�JJJ�RRR�TTT�SSS�>>>�BBB�HHH�PPP�SSS�WWW�ZZZ�]]]�```�ddd�hhh�```�VVV�VVV�WWW�VVV�VVV�VVV�WWW�kkk�ooo�ooo�nnn�ppp�ooo�ggg�hhh�hhh�ggg�hhh�hhh�ggg�ggg�mmm�nnn�ppp�rrr�xxx�zzz�����������������������������x�x�v�v�s�t�p�q�o�p�o�p�{�{�����uuu�sss�����������������pppY   /   $                     ��� ��� ��� ��� ���                 ��                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���+���Y���`zzz�uuu��   �!!!�---�888�;;;�LLL�TTT�WWW�UUU�>>>�AAA�GGG�QQQ�TTT�XXX�[[[�___�aaa�fff�iii�aaa�XXX�XXX�WWW�VVV�WWW�WWW�XXX�mmm�ppp�ppp�qqq�rrr�qqq�hhh�iii�iii�iii�iii�iii�jjj�iii�mmm�qqq�ppp�sss�zzz�zzz�����������������������������~�~�|�|�w�w�w�x�y�z�~�~�����uuu�ttt�ttt�����������������pppY   /   $                     ��� ��� ��� ��� ��� ��� ���                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���+���Y���`����|||��   �"""�...�888�;;;�NNN�VVV�XXX�WWW�???�CCC�III�QQQ�UUU�YYY�\\\�___�bbb�fff�jjj�ccc�XXX�YYY�XXX�XXX�XXX�YYY�YYY�ooo�rrr�sss�sss�rrr�rrr�jjj�jjj�jjj�kkk�kkk�lll�kkk�kkk�ooo�rrr�qqq�ttt�{{{�}}}���������������������������������������|�|���������xxx�vvv�ttt�uuu�����������������pppY   /   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���+���Y���_����|||��!!!�###�///�:::�<<<�PPP�YYY�ZZZ�XXX�???�CCC�HHH�RRR�VVV�YYY�\\\�```�ddd�ggg�kkk�aaa�YYY�ZZZ�XXX�YYY�YYY�YYY�ZZZ�ppp�sss�ttt�ttt�vvv�ttt�kkk�lll�lll�mmm�lll�mmm�mmm�mmm�qqq�rrr�ttt�uuu�|||�~~~�����������������������������������������������������www�www�vvv�vvv�����������������pppY   /   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���+���X���_����}}}��!!!�###�///�;;;�>>>�QQQ�ZZZ�\\\�ZZZ�>>>�CCC�III�SSS�WWW�[[[�^^^�```�ddd�iii�kkk�ccc�ZZZ�[[[�ZZZ�YYY�[[[�[[[�ZZZ�qqq�uuu�vvv�vvv�www�vvv�nnn�mmm�mmm�nnn�nnn�nnn�mmm�mmm�rrr�uuu�ttt�www�~~~���������������������������������������������������������xxx�xxx�www�www�zzz�|||���������oooY   /   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���*���X���_����}}}��"""�###�000�;;;�>>>�RRR�\\\�^^^�\\\�???�CCC�JJJ�SSS�XXX�[[[�___�bbb�eee�iii�mmm�ddd�ZZZ�\\\�[[[�YYY�ZZZ�[[[�[[[�ttt�vvv�xxx�xxx�xxx�xxx�nnn�nnn�ooo�ooo�ppp�ppp�ooo�ooo�uuu�vvv�uuu�xxx�������������������������������������������������������������zzz�yyy�www�xxx�sss�uuu���������oooY   /   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���*���W���^����}}}��!!!�$$$�111�===�@@@�TTT�___�```�]]]�???�CCC�JJJ�TTT�XXX�\\\�___�ccc�fff�jjj�nnn�ddd�ZZZ�\\\�[[[�\\\�[[[�\\\�]]]�ttt�zzz�zzz�yyy�zzz�{{{�ppp�ooo�ooo�ppp�qqq�qqq�qqq�qqq�vvv�www�www�zzz�������������������������������������������������������������zzz�zzz�xxx�xxx�ttt�nnn���������oooY   /   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���*���W���^����}}}�   �"""�$$$�222�>>>�AAA�VVV�aaa�bbb�```�@@@�DDD�JJJ�UUU�YYY�]]]�___�ccc�ggg�kkk�ooo�ddd�ZZZ�]]]�\\\�[[[�\\\�\\\�]]]�vvv�{{{�{{{�{{{�{{{�{{{�qqq�qqq�rrr�rrr�rrr�sss�sss�sss�yyy�yyy�xxx�{{{�������������������������������������������������������������zzz�zzz�zzz�zzz�{{{�uuu���������oooY   /   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���*���W���^����}}}�   �"""�$$$�333�???�BBB�WWW�bbb�eee�bbb�@@@�DDD�KKK�UUU�ZZZ�]]]�```�eee�hhh�kkk�ooo�eee�ZZZ�]]]�]]]�\\\�]]]�\\\�]]]�www�|||�|||�}}}�}}}�~~~�sss�sss�sss�ttt�ttt�uuu�ttt�ttt�zzz�{{{�zzz�}}}�������������������������������������������������������������{{{�|||�zzz�{{{�����}}}���������oooY   /   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���)���W���^����}}}�   �"""�%%%�333�@@@�CCC�XXX�eee�ggg�ccc�AAA�EEE�KKK�VVV�[[[�___�aaa�eee�iii�mmm�ooo�eee�ZZZ�]]]�]]]�^^^�]]]�^^^�^^^�yyy�~~~�~~~�������ttt�uuu�ttt�uuu�uuu�uuu�ttt�vvv�zzz�|||�{{{�~~~�������������������������������������������������������������}}}�|||�{{{�{{{�����������������oooW   /   $                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���)���V���\����}}}�!!!�"""�$$$�555�BBB�DDD�[[[�hhh�iii�ddd�AAA�DDD�KKK�VVV�ZZZ�___�aaa�eee�iii�mmm�ppp�ggg�YYY�]]]�^^^�]]]�]]]�___�___�{{{������������������vvv�vvv�vvv�www�vvv�www�vvv�www�|||�~~~�|||�����������������������������������������������������������������}}}�}}}�}}}�{{{�����������������oooW   .   #                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 	���)���U���\����}}}�!!!�###�%%%�555�CCC�EEE�\\\�hhh�kkk�fff�AAA�EEE�LLL�WWW�\\\�___�bbb�fff�jjj�nnn�qqq�fff�YYY�]]]�^^^�^^^�^^^�___�aaa�}}}���������������������vvv�www�vvv�www�www�www�xxx�xxx������}}}�����������������������������������������������������������������~~~�}}}�|||�|||�����������������oooV   -   "                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 ���(���T���Z����}}}�"""�$$$�%%%�666�DDD�FFF�^^^�kkk�nnn�hhh�@@@�EEE�LLL�XXX�]]]�___�ccc�fff�kkk�nnn�rrr�fff�ZZZ�\\\�^^^�___�```�```�```�~~~���������������������xxx�yyy�xxx�xxx�yyy�zzz�zzz�zzz���������������������������������������������������������������������������~~~�~~~�~~~�����������������qqqT   ,   !         
            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 ���'���S���Y����~~~�###�$$$�%%%�777�EEE�GGG�___�nnn�ppp�jjj�@@@�DDD�LLL�YYY�]]]�```�ddd�ggg�kkk�nnn�sss�fff�YYY�^^^�^^^�___�aaa�```�aaa����������������������zzz�zzz�zzz�{{{�zzz�zzz�{{{�zzz�������������������������������������������������������������������������������~~~�}}}�����������������uuuR   )            	             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 ���'���R���X����}}}�###�%%%�&&&�888�FFF�III�aaa�ppp�rrr�mmm�@@@�FFF�MMM�XXX�^^^�aaa�ddd�hhh�lll�ppp�sss�fff�ZZZ�]]]�^^^�___�```�```�bbb�������������������������{{{�|||�{{{�|||�|||�|||�|||�|||������������������������������������������������������������������������������~~~�~~~�}}}�����������������yyyO   &            	             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                         ��� ��� ��� ��� ��� ���                 ���%���P���U����~~~�$$$�&&&�&&&�888�HHH�KKK�ccc�sss�ttt�ooo�AAA�FFF�MMM�YYY�^^^�aaa�ddd�hhh�lll�qqq�sss�ggg�YYY�]]]�^^^�```�aaa�bbb�bbb�������������������������|||�}}}�}}}�}}}�}}}�}}}�}}}�~~~�����������������������������������������������������������������������������~~~�}}}�|||�{{{��������������������K   #                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                 ��� ��� ��� ���                  ���$���N���S����~~~�$$$�&&&�'''�999�JJJ�LLL�ddd�ttt�vvv�qqq�AAA�EEE�NNN�ZZZ�^^^�bbb�eee�iii�mmm�ppp�uuu�ggg�YYY�^^^�^^^�___�aaa�bbb�bbb�������������������������}}}�}}}�~~~�~~~�~~~�����������������������������������������������������������������������������������}}}�{{{�{{{�{{{�������������������F            
                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                          ��� ���                  ���"���L���P��������&&&�'''�(((�:::�KKK�NNN�ggg�www�yyy�rrr�AAA�FFF�MMM�[[[�___�bbb�fff�jjj�nnn�qqq�vvv�iii�YYY�]]]�^^^�```�aaa�ccc�ccc����������������������������������������������������������������������������������������������������������������������������}}}�{{{�{{{�zzz���������������z���A            	                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                          ��� ���              ���!���J���N��������CCC�'''�(((�<<<�LLL�OOO�iii�yyy�|||�ttt�AAA�FFF�MMM�ZZZ�___�bbb�fff�jjj�ooo�rrr�uuu�iii�XXX�\\\�]]]�___�bbb�ddd�ccc����������������������������������������������������������������������������������������������������������������������������������{{{�zzz�yyy����������������y���v���;         
                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                             ������H���L���ć���uuu�AAA�***�===�NNN�PPP�jjj�|||�~~~�www�AAA�EEE�NNN�[[[�```�ccc�ggg�kkk�nnn�rrr�xxx�iii�YYY�]]]�]]]�___�bbb�ccc�ddd�������������������������������������������������������������������������������������������������������������������������������������zzz�zzz��������������������t���q���.                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                            ������H���J���N������������������������������������������������������������������������������������������������������������������������������������������������������ttt�iii�eee�ppp�|||����������������������������������������������������������������������������������������������������s���o���mddd                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                      	   
      
   	                                            ���-���H���K���O���ǌ��򋋋���������������������������������������������������������������������������������������������������������������������������������������������vvv�iii�]]]�ggg�ttt������������������������������������������������������������������������������������������������r���n���k���F   
                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                	                        
                                    iii���5���J���M���O���T���[����а�׿�����鉉�������������������������������������������������ٝ��|���u���o���i���e���a���^���]���\���\���[���[���\���\���]���]���^���^���^���_���_���`���b���c���g���k�����������������������������������������������������������������������z���u���p���m���j���L\\\                          ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                  ������/���;¿�D���r�ͦ�ڷ|�ɥg}����{{{�����������������������������������������}}}�����i���a���Y���R���L���G���D���A���@���?���@���@���@���@���@���A���A���A���A���B���B���D���E���G���K���O�����������������������������������������������������������v���o���g���`���Y���R���B���(   	                          ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���             
���+�γ�F<2                           	                                 	      OD9�ĬW翄�י:s�v _�qbqme�\\\�������������������������������������kkk�\\\�___�   A   6   +   !               	                                          	         bbb�\\\�������������������������������������___�\\\�999|   H   =   2   '            
                          ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���          	   �д��Ѱ��̰�7/'                            	                           	   
   SSG�ȳ^�Ŋ��=z�} d�v d�tfrmd�\\\�������������������������������������kkk�\\\�``^�   @   5   *                                                                	      bbb�\\\�������������������������������������___�\\\�999|   G   <   1   %                                    ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���          	�¦d�Ҳ������ά��Ȯ�0)"%                            	                     	      [OO�̴h�Ǝ��?�Ձ k�| i�x h�sksmd�\\\�������������������������������������kkk�\\\�a`^� C   4   )                                                                     bbb�\\\�������������������������������������___�\\\�999{   F   ;   0   $                             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       �� �ѳ��Ě��v���d��ϭ��Ǭ�*$*   #   !                        	         	   
      ^SI�Ͷp�Ǒ��A�ۂ r� o�} n�x m�vosmc�\\\�������������������������������������kkk�\\\�ca]�! F 8   )            
                                                           bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   $                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       �ǫv�ѳ���7��q ��r ���e��έ��ū�("-   %   #                                    aWM�εx�Ȕ��C�߁ zۂ x� t�z s�x r�vtsmc�\\\�������������������������������������kkk�\\\�db]�1# J' ; .                                              ��� ���                       bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       	�̮��ѱ��r��p ��q ��q ���d��Ϭ��é�&!/   '   #                               `OF�͵��ɖ��C�� ��� �� |� {�{ x�v v�wytmc�\\\�������������������������������������kkk�\\\�ec\�>* N8( @. 2# $                                       ��� ��� ���                       bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       	�ή������n ��o ��p ��p ��q ���c��Ϭ�����%1   (   $   !                     ZRJ�δ��ș��F�� �� ��� �� ��| �| }�w |�u}unb�\\\�������������������������������������kkk�\\\�gc\�H2 QG1 DB/ 6:& (-$                                         ��� ���                       bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �|c�а���n��m ��m ��o ��o ��p ��p ���c��ϭ��¨�$2   (   %   !               UN@$�˳��ʜ��F�� ��~ �� ��} ��~ ��} ��z ��y ��w�unb�\\\�������������������������������������kkk�\\\�hd\�S8 VQ9 HR8 ;O8 -G0  ;/                                     ��� ���                       bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ͦ�(�ͮ���Y��l ��l ��m ��n ��o ��p ��p ���c��ή�����$2   )   &   #   !      RE?)�̲��ɞ��G��} ��} ��} ��} ��~ ��| ��| ��{ ��w ��y�vnb�\\\�������������������������������������kkk�\\\�hd[�^? Z^@ L^B >bC 2aF %Z< L= FFF+++                           ��� ���                       bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    Ȝ�)�̬���W��k ��k ��l ��m ��n ��o ��o ��p ���c��Ϯ�����#3   *   (   %   #MB7.�ɱ��ʠ��H��{ ��{ ��| ��| ��| ��| ��} ��{ ��z ��y ��w�vna�\\\�������������������������������������kkk�\\\�je[�fE ]iF PlI BoM 5sO *wU pJ ��[���                            ��� ���                       bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    Ȝ�)�˪���V��i ��k ��k ��l ��m ��n ��o ��o ��p ���b��έ��§�#4   ,   *E;64�ȭ��ʢ���I��z ��z ��z ��z ��{ ��{ ��{ ��{ ��{ ��y ��x ��y�wna�\\\�������������������������������������kkk�\\\�ke[�oJ `qM SwP F|T 9�Y .�_ #�k
īr���                        ��� ��� ���                       bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    Ȝ�)�ʩ���U��h ��i ��j ��k ��l ��l ��n ��n ��o ��p ���b��Ϯ�����"5B90:�Ƭ��ͥ���J��x ��y ��y ��y ��z ��z ��{ ��{ ��z ��z ��z ��w ��y�xna�\\\�������������������������������������kkk�\\\�mfY�vM c{R W�V J�[ >�b 1�j &Ȣ\/Ҽ�#��u                        ��� ��� ���                       bbb�\\\�������������������������������������___�\\\�999{   F   ;   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    Ȝ�)�ȧ���T��g ��h ��i ��j ��k ��l ��l ��n ��n ��o ��p ���b��ϯ��¨��Ƭ��ͩ���K��v ��v ��x ��x ��y ��y ��y ��y ��z ��z ��z ��y ��x ��w�xn`�\\\�������������������������������������kkk�\\\�nfY�~R g�U Z�[ O�b A�h 6ȤX@Ѻ�7���                                                           bbb�\\\�������������������������������������___�\\\�:::{   F   :   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ę{*�ǥ���S��f ��g ��h ��i ��j ��k ��l ��l ��n ��n ��o ��p ���b��Я��Ϋ���K��s ��u ��u ��u ��w ��x ��y ��y ��y ��y ��z ��y ��x ��w ��y�yn`�\\\�������������������������������������kkk�\\\�ngYՅU l�Y _�] R�e FŠSSҶ�I���$                                                         bbb�\\\�������������������������������������___�\\\�:::{   F   :   /   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ę{*�ţ���S��f ��f ��g ��h ��i ��j ��k ��k ��l ��n ��n ��o ��p ���b���M��r ��s ��s ��u ��u ��u ��w ��w ��x ��y ��x ��x ��y ��x ��w ��{�zo_�\\\�������������������������������������kkk�\\\�pgX֊W o�\ d�a WRf̳�\���1      	                                                	      bbb�\\\�������������������������������������___�\\\�:::{   E   :   .   #                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ē{*�ġ���R��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��n ��n ��o ��p ��p ��r ��r ��s ��s ��u ��u ��u ��w ��w ��x ��x ��x ��x ��x ��z��z
�zo_�\\\�������������������������������������kkk�\\\�qhX؏Z t�^h��Ryɰ�p���?                                                      	         bbb�\\\�������������������������������������___�\\\�:::{   D   9   -   "         
             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ē{*�à���Q��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��m ��n ��o ��p ��p ��q ��r ��s ��s ��u ��u ��u ��w ��w ��x ��x ��x ��{��{��z	�{o_�\\\�������������������������������������kkk�\\\�rhWڕ^z��Q�Ū�����N                	                                 	   
            bbb�\\\�������������������������������������___�\\\�:::z   D   8   ,   !         
             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ē{*������P��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��m ��n ��o ��p ��p ��q ��r ��s ��s ��u ��u ��u ��w ��w ��x ��{��z��z��z	�{n_�\\\�������������������������������������mmm�]]]�tiW���Q�è����y_,   #                                                                bbb�\\\�������������������������������������___�\\\�;;;y   B   7   +   !         	             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��r*������O��b ��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��m ��n ��o ��p ��p ��q ��r ��s ��s ��u ��u ��u ��w ��{��|��z��z��y�{o_�]]]�������������������������������������ppp�```��wi�ĩ���~so:   1   )   "                                                         !   'aaa�\\\�������������������������������������___�\\\�;;;w   A   6   *            	             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��r*������N��a ��b ��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��m ��n ��o ��p ��p ��q ��r ��s ��s ��u ��u��y��{	��{��z��z��z��q]�___�������������������������������������yyy�ccc�}xsw�K   ?   7   0   *   %   "                                             !   $   )   /```�\\\�������������������������������������]]]�\\\�%%%a   ?   3   (            	             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��r*�����M��` ��a ��b ��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��m ��n ��o ��p ��p ��q ��r ��s ��s��y	��z
��y	��{��y��z��{��wV�bbb�|||�������������������������������������fff�onn�!!!\SI@   9   3   /   ,   )   (   '   &   &   &   &   &   &   &   &   '   (   )   +   .   2   7]]]�\\\�������������������������������������\\\�]]]�   G   <   1   &                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��r*�����L��` ��` ��a ��b ��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��m ��n ��o ��p ��p ��q ��r��x
��z��z
��z	��y��y��{	��}��~L�ddd�sss�������������������������������������hhh�iii�>>>x"""[SK   B   =   9   6   4   3   2   1   1   1   1   1   1   1   1   2   3   4   6   9   =]]]�\\\�```�������������������������������������\\\�^^^�   D   9   .   #                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��l*������K��_ ��` ��` ��a ��b ��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��m ��n ��o ��p ��r��v��x��z��x
��z	��y��z
��~���̓3�fff�kkk�������������������������������������vvv�iii�mmm�'''b!!!\UN   G   D   A   @   ?   >   =   =   =   =   =   =   =   =   >   >   ?   A   D111e___�\\\�}}}�������������������������������������\\\�___�   @   6   *             
            ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��l*�����K��^ ��_ ��` ��` ��a ��b ��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��m ��n ��p��v
��x��x��x��x
��x	��z	��|��~�����nnm�kkk�����������������������������������������mmm�jjj�mmm�XXX�]XQ   M   L   J   I   H   H   H   H   H   H   H   H   H   H   I   JS\\\�^^^�\\\�fff�������������������������������������nnn�\\\�aaa�   <   1   '            	             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��l*�����J��] ��^ ��_ ��` ��` ��a ��b ��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��k ��l ��o��u��v��w��w��x��w
��x��y��~������ Ƅyn�mmm���������������������������������������������ppp�iii�hhh�fff�fff�ccc�___�```�```�```�```�```�```�```�```�```�```�```�```�```�```�___�]]]�\\\�\\\�hhh�����������������������������������������___�\\\�SSS�   7   ,   #                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��j+�����I��\ ��] ��^ ��_ ��` ��` ��a ��b ��c ��d ��e ��f ��f ��g ��h ��i ��j ��k ��l��s��v��v��v��v��w
��v	��w
��z��}������ȵ�Y�ooo�vvv����������������������������������������������mmm�fff�ddd�```�]]]�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�ddd����������������������������������������������\\\�^^^�   ;   1   (            
                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��j+�����H��[ ��\ ��] ��^ ��_ ��` ��` ��a ��b ��c ��d ��e ��f ��f ��g ��h ��i ��k��r��s��t��u��v��u��v
��u
��x��z��~������!��*�xvt�sss�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ddd�\\\�bbb�   5   ,   "                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��d+�����G��Z ��[ ��\ ��] ��^ ��_ ��` ��` ��a ��b ��c ��d ��e ��f ��f ��g ��i��p��s��s��s��s��u��u��u��u
��x��z��~�������$��+ΰ�d�ttt�~~~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������\\\�^^^�E   /   %            
                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��d+�����F��Y ��Z ��[ ��\ ��] ��^ ��_ ��` ��` ��a ��b ��c ��d ��e ��f ��g��o��q��r��r��s��r��s��t��u��t
��w��z��~�������%���*��4Ђ�~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������```�\\\�aaa�   0   (                               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��d+�����E��Y ��Y ��Z ��[ ��\ ��] ��^ ��_ ��` ��` ��a ��b ��c ��d ��f��n��p��p��q��q��r��r��r��r��t��s
��v��z��}���� ��%��,�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ddd�\\\�```�4   )   !            	                ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��d+�����D��X ��Y ��Y ��Z ��[ ��\ ��] ��^ ��_ ��` ��` ��a ��b ��d��m��p��p��p��p��p��q��q��r��q��r��s
��u��y��|���� ��'������׽��ʷ�������������������������������������������������������������������������������������������������������������������������������������������������������������������������iii�\\\�___�000K   )   !            
                    ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��d+�����D��W ��X ��Y ��Y ��Z ��[ ��\ ��] ��^ ��_ ��` ��` ��b��l��n��o��o��p��o��p��p��q��q��r��q
��r
��u��x��{�����������׽��ȳ���X���e���ݘ�����������������������������������������������������������������������������������������������������������������������������������������������������������ccc�\\\�^^^�TTTs   (   !                               ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ��^+�����C��V ��W ��X ��Y ��Y ��Z ��[ ��\ ��] ��^ ��_ ��a��j��m��n��n��n��o��o��o��o��p��p��q��q
��q	��s��x��y��}������y��׾��͵˄}X���]���k���Ӗ�����������������������������������������������������������������������������������������������������������������������������������������������|||�___�\\\�___�QQQm   %                                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �~`*�����B��U ��V ��W ��X ��Y ��Y ��Z ��[ ��\ ��] ��_��j��m��l��m��m��n��n��n��o��n��o��o��p��p
��q
��q��u��x��{��~��� ���z��ٿ��̷͉��Y���_���h��������������������������������������������������������������������������������������������������������������������������������������������ccc�\\\�\\\�```�555C   "                                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �~`*�����A��T ��U ��V ��W ��X ��Y ��Y ��Z ��[ ��]��i��l��l��l��l��l��m��m��n��n��n��n��n��o��o
��p
��q
��s��v��z��|�����"���|��ٿ��η̇��X���Y���^���z����zzz�uuu�sss�zzz�������������������������������������������������������������������������������������������������}}}�lll�]]]�\\\�\\\�^^^�ddd�%                  
                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    āb*��~��@��S ��T ��U ��V ��W ��X ��Y ��Y ��[��g��k��k��k��l��l��k��l��l��m��m��n��n��m��n��n��o
��o	��r��t��w��z��}�����!���{��ؾ��η̇�U}}}P���O���O���|||�sss�ooo�mmm�jjj�hhh�eee�ccc�```�]]]�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�___�eee�###*                     	                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    ͆`(��|��~?��S ��S ��T ��U ��V ��W ��X ��Z��f��i��j��j��j��k��k��l��k��k��l��l��m��m��m��m��m��n
��n	��p
��r��v��w��{��~������ ���{��ؽ��ͷ́||QyyyJ{{{H|||F~~~D���H����xxx�qqq�kkk�ggg�aaa�___�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�\\\�]]]�^^^�```�aaa�eee�YYYc                        	                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���    �sS��z��F��R ��S ��S ��T ��U ��V ��X��e��i��i��i��i��j��j��j��k��k��k��k��k��l��l��m��m��m��m
��m	��n��p
��s��v��w��z��}��������x��׽��ε�}wwLpppBppp@sss<uuu9rrr5rrr1sss.ppp*ggg']]]-ZZZ4WWW3ZZZ4ZZZ4ZZZ4ZZZ4WWW3WWW3SSS2PPP1III/AAA.<<<-888,888,888,                                 	                             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ��w��]��Q ��R ��S ��S ��T ��V��d��h��h��i��h��h��i��i��i��j��j��k��j��k��k��k��l��l��m��l
��m	��m��n��p��s��v��v��z��}��~�����x��ֺ��̵�yrrDiii:hhh6jjj2hhh,ggg'ddd$ZZZFFF...                                          	                                   ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ��v���s��Q��Q ��R ��S ��T��c��g��g��g��h��h��h��h��h��i��i��i��j��j��j��j��j��k��k��l��l
��l
��l	��m��n��p
��r��u��w��y��z��}��}���v��չ��Ͳ�skk;^^^1bbb,]]]']]]!TTTGGG---            
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   	   	   	                                             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       ��r���v��^��P ��Q ��S��c��f��f��f��g��g��g��h��g��g��h��h��i��i��i��j��i��j��j��j��k��k
��l
��k	��l��l��n��o	��r
��s��v��w��y��y��{���s��Է��˱�pff1QQQ&OOO MMM>>>000      	                                                                                                      ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���       �j<��u��R��O ��Q��a��e��f��e��f��f��f��g��g��g��g��g��g��h��h��h��i��i��i��i��j��j��j��k
��k	��k��k��l��l��n��o��r	��s��v��v��x��x���p��ӵ��̰�ic\&<<<444"""                                                                                                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���          ��r���t��m,��`��d��e��e��e��e��e��e��f��f��f��g��f��g��g��g��h��h��h��i��h��i��i��j��j
��j	��k��j��k��k��l��n��n��o��q��s��t��u��v���o��Ҵ��̯�`WN                                                                                                       ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���          �gE��q���x��l*��d��d��d��e��e��d��e��e��e��f��f��f��f��f��f��g��g��h��h��h��h��h��i��i
��j	��j��j��j��j��k��k��m��m��n��n��p��q��s��s���j��Ѳ��ͮ�m`R   	                                                                                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���              �i=��s���|�فG��c��c��d��d��d��d��d��d��e��e��e��f��e��f��f��f��g��g��g��h��g��h��h
��i	��i��j��j��j��j��j��k��l��m��m��n ��o ��q ��r �����ɤ��в��ͯ�                          ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 �k4��p���}��i��v8��g#��c��c��d��c��d��d��d��e��e��e��e��e��f��f��f��g��g��g��g��g
��h	��h	��i��i��j��i��j��j��j��l��l��m ��n��~���X��˩��έ��ʬ��zk                       ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                 �^F��p���w����������x��c��^��_��^��_��`��`��_��`��`��a��a��a��b���b���b���c���c���d���c���d���d���d���e���e���f���f���g���g���i�����Ġ��ɨ��ʪ��ʨ�巜8                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                     �f*��og��r���w���x���{���|���~�����������������������������������������������������������������������������������������������à��Ţ��š��ģ��¡��M`@@                             ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                                                                                     ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��������������������������������������������������������������������������������������������������������������������������    �����������    �����������    �����������    �����������     �����������     ����������     ����������     ?����������     ?����������     ?�����������    ?�����������    ?�����������    ?�����������    ?�����������    ?�����������    ?�����������    ?�����������    ?�����������    ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����           ?����         ` ?����         � ?����        � ?����        � ?����        � ?����        � ?����        ��?����        ������        ������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        �������        ?�������        �������        �������        �������        ��������       ��������� ��� ��������  ��� ��������� ��� ���������� ��� ���������� ��� ��������� ��� ������?��� ��� ��������� ��� �������� ��� �������   ��� �������   ��� �������   ��� ������ �   ��� ������ `   ��� ������     ��� ������     ��� ������     ��� ������     ��� ������     O��� ������     ��� ������     ?��� ������     ?��� ������     ��� ������     ��� ������     ?��� ������     ��  ������          ������         ������         ������         ������         ������         ������         ������        ������   �    ?������   �    ������    �    �������    |   �������    ?   �������    �����������    �����������    �����������    �����������    �����������     �����������     ����������     ?����������     ����������    ������������   ��������������������������Transparent	  TLabelLabel3LeftHTop/Width[HeightAnchorsakLeftakBottom Caption   Copyright för vissa delar:  TLabelRegistrationLabelLeftHTop� WidthHeightAnchorsakLeftakBottom CaptionThis product is licensed to:  TStaticTextHomepageLabelLeftHTopHWidth� HeightCaptionhttp://XXXXXXwinscp.net/TabOrderTabStop	  TStaticTextForumUrlLabelLeftHToptWidth� HeightCaptionhttp://XXXXwinscp.net/forum/TabOrderTabStop	  TStaticTextTranslatorUrlLabelLeftHTop� Width� HeightCaptionhttp://XXXXwinscp.net/forum/TabOrderTabStop	  
TScrollBoxThirdPartyBoxLeftHTopAWidth2HeightyHorzScrollBar.Range!HorzScrollBar.VisibleVertScrollBar.Range�VertScrollBar.Smooth	VertScrollBar.Tracking	AnchorsakLeftakRightakBottom 
AutoScrollTabOrder
DesignSizeu  TLabelLabel7LeftTopWidth� Height)AnchorsakLeftakTopakRight AutoSizeCaptionW   Licensavtalen för följande program (bibliotek) är del av applikationens licensavtal.WordWrap	  TLabelPuttyVersionLabelLeftTop0Width� HeightCaption#SSH and SCP code based on PuTTY xxx  TLabelPuttyCopyrightLabelLeftTop@Width� HeightCaption   Copyright © xxx Simon Tatham  TLabelLabel8LeftTopmWidth� HeightCaption'Filemanager Toolset library Version 2.6  TLabelLabel10LeftTop}Width� HeightCaption   Copyright © 1999 Ingo Eckel  TLabelLabel1LeftTop� WidthzHeightCaptionToolbar2000 library 2.1.6  TLabelLabel2LeftTopWidth� HeightCaption%   Copyright © 1998-2005 Jordan Russell  TLabelLabel5LeftTop5WidthFHeightCaptionTBX library 2.1  TLabelLabel6LeftTopEWidth� HeightCaption&   Copyright © 2001-2005 Alex A. Denisov  TLabelFileZillaVersionLabelLeftTop� Width� HeightCaptionFTP code based on Filezilla xxx  TLabelFileZillaCopyrightLabelLeftTop� Width� HeightCaption   Copyright © xxx Tim Kosse  TLabelOpenSSLVersionLabelLeftTop� WidthHeightAutoSizeCaptioncThis product includes software developed by the OpenSSL Project for use in the OpenSSL Toolkit xxx.WordWrap	  TLabelOpenSSLCopyrightLabelLeftTop� Width� HeightCaption%   Copyright © xxxx The OpenSSL Project  TStaticTextPuttyLicenseLabelTagLeftTopPWidthIHeightCaptionVisa licensTabOrder TabStop	OnClickPuttyLicenseLabelClick  TStaticTextPuttyHomepageLabelLeftTop`WidthHeightCaption5http://XXXwww.chiark.greenend.org.uk/~sgtatham/putty/TabOrderTabStop	  TStaticTextToolbar2000HomepageLabelLeftTopWidth� HeightCaption$http://www.jrsoftware.org/tb2kdl.phpTabOrderTabStop	  TStaticTextTBXHomepageLabelLeftTopUWidth� HeightCaption!https://github.com/plashenkov/TBXTabOrderTabStop	  TStaticTextFileZillaHomepageLabelLeftTop� Width� HeightCaption$http://XXXfilezilla.sourceforge.net/TabOrderTabStop	  TStaticTextOpenSSLHomepageLabelLeftTop� WidthvHeightCaptionhttp://XXX.openssl.org/TabOrderTabStop	   TButtonOKButtonLeft� Top�WidthKHeightAnchorsakRightakBottom Cancel	CaptionOKDefault	ModalResultTabOrder OnMouseDownOKButtonMouseDown  TButtonLicenseButtonLeftHTop�WidthKHeightAnchorsakLeftakBottom Caption
&Licens...TabOrderOnClickLicenseButtonClick  TButton
HelpButtonLeft/Top�WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  
TScrollBoxRegistrationBoxLeftHTop� Width2HeightYHorzScrollBar.VisibleVertScrollBar.Smooth	VertScrollBar.Tracking	AnchorsakLeftakRightakBottom TabOrder
DesignSize.U  TLabelRegistrationSubjectLabelLeftTopWidthHeightAAnchorsakLeftakTopakRight AutoSizeCaptionSomeone
Somewhere, some cityWordWrap	  TLabelRegistrationLicensesLabelLeftTop+WidthjHeightCaptionNumber of Licenses: X  TStaticTextRegistrationProductIdLabelLeftTopAWidth� HeightCaptionProduct ID: xxxx-xxxx-xxxxxTabOrder OnClickRegistrationProductIdLabelClick      TPF0TAuthenticateFormAuthenticateFormLeft0TopqHelpType	htKeywordHelpKeywordui_authenticateBorderIconsbiSystemMenu BorderStylebsDialogCaptionAuthenticateFormClientHeightgClientWidthwColor	clBtnFaceConstraints.MinHeight� Constraints.MinWidth
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnResize
FormResizeOnShowFormShowPixelsPerInch`
TextHeight 	TListViewLogViewLeft Top WidthwHeight,AlignalClientColumnsWidthd  DoubleBuffered	ReadOnly		RowSelect	ParentDoubleBufferedShowColumnHeadersTabOrder 	ViewStylevsReport  TPanelPasswordPanelLeft Top,WidthwHeight� AlignalBottomAutoSize	
BevelOuterbvNoneTabOrderVisible TPanelPromptEditPanelLeft Top WidthwHeight� AlignalTop
BevelOuterbvNoneTabOrder 
DesignSizew�   TLabelInstructionsLabelLeftTopWidthhHeight'AnchorsakLeftakTopakRight AutoSizeCaption�Instructions for authentication. Please fill in your credentials carefully. Enter all required information, including your session username and session password.XFocusControlPromptEdit1WordWrap	  TLabelPromptLabel1LeftTop8WidthhHeightAnchorsakLeftakTopakRight AutoSizeCaption&UsernameX:FocusControlPromptEdit1WordWrap	  TLabelPromptLabel2LeftTopeWidthhHeightAnchorsakLeftakTopakRight AutoSizeCaption&PasswordX:FocusControlPromptEdit2WordWrap	  TPasswordEditPromptEdit1LeftTopIWidthiHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder   TPasswordEditPromptEdit2LeftTopvWidthiHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder   TPanelSavePasswordPanelLeft Top� WidthwHeightAlignalTop
BevelOuterbvNoneTabOrder 	TCheckBoxSavePasswordCheckLeftTopWidthHeightCaption   &Ändra lösenord till det härChecked	State	cbCheckedTabOrder    TPanelButtonsPanelLeft Top� WidthwHeight,AlignalTop
BevelOuterbvNoneTabOrder
DesignSizew,  TButtonPasswordOKButtonLeftvTopWidthKHeightAnchorsakTopakRight CaptionOKModalResultTabOrder   TButtonPasswordCancelButtonLeft� TopWidthKHeightAnchorsakTopakRight CaptionAvbrytModalResultTabOrder  TButtonPasswordHelpButtonLeft&TopWidthKHeightAnchorsakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick   TPanelSessionRememberPasswordPanelLeft Top� WidthwHeightAlignalTop
BevelOuterbvNoneTabOrder 	TCheckBoxSessionRememberPasswordCheckLeftTopWidthHeightCaption.   &Kom ihåg lösenordet för den här sessionenChecked	State	cbCheckedTabOrder     TPanelBannerPanelLeft TopWidthwHeightRAlignalBottom
BevelOuterbvNoneTabOrderVisible
DesignSizewR  TMemo
BannerMemoLeftTopWidthhHeight"AnchorsakLeftakTopakRightakBottom Color	clBtnFaceReadOnly	
ScrollBars
ssVerticalTabOrder WantReturns  	TCheckBoxNeverShowAgainCheckLeftTop5Width� HeightAnchorsakLeftakRightakBottom Caption&   &Visa aldrig det här meddelandet igenTabOrder  TButtonBannerCloseButtonLeft� Top/WidthKHeightAnchorsakRightakBottom Caption	   FortsättModalResultTabOrder  TButtonBannerHelpButtonLeft$Top/WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick     TPF0TCleanupDialogCleanupDialogLeftdTop� HelpType	htKeywordHelpKeyword
ui_cleanupBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionRensa applikationsdataClientHeight+ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnShowFormShow
DesignSize�+ PixelsPerInch`
TextHeight TLabelLabel1LeftTopWidth�HeightaAnchorsakLeftakTopakRight AutoSizeCaption8  Följande lista innehåller all data som det här programmet lagrar på den här datorn. Välj det som du vill ska tas bort.

Om ytterligare instanser av programmet är igång, var god avsluta dem innan nedanstående data tas bort.

Notera att en del av dessa data kommer att återskapas vid nästa uppstart.WordWrap	  TButtonOKButtonLeft� TopWidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeftITopWidthKHeightAnchorsakRightakBottom Cancel	Caption   StängModalResultTabOrder  	TListViewDataListViewLeftTophWidth�Height� AnchorsakLeftakTopakRightakBottom 
Checkboxes	ColumnsCaptionDataTagWidth�  CaptionPlatsWidth�  ColumnClickDoubleBuffered	HideSelectionReadOnly		RowSelect	ParentDoubleBufferedParentShowHintShowHint	TabOrder 	ViewStylevsReport	OnInfoTipDataListViewInfoTipOnKeyUpDataListViewKeyUpOnMouseDownDataListViewMouseDown  TButtonCheckAllButtonLeftTop
WidthlHeightAnchorsakLeftakBottom CaptionMarkera &allaTabOrderOnClickCheckAllButtonClick  TButton
HelpButtonLeft�TopWidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick   TPF0TConsoleDialogConsoleDialogLeft]Top� HelpType	htKeywordHelpKeyword
ui_consoleBorderIconsbiSystemMenu
biMaximizebiHelp CaptionKonsolClientHeight�ClientWidth'Color	clBtnFaceConstraints.MinHeight� Constraints.MinWidth�
ParentFont		Icon.Data
~           h     (                 @                                                                                  '!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�(!�'!�'!�/'"�/'"�/'"�/'"�/'"�/'"�/'"�/'"�/'"�/'"�/'"�/'"�/'"�/'"�'!�'!�SJE�����rje�6-'�6-'�6-'�6-'�6-'�6-'�6-'�6-'�6-'�6-'�6-'�'!�'!�=3,�d[U���������PF@�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�=3,�'!�'!�D91�D91�SHA���������D91�D91�D91�D91�D91�D91�D91�D91�D91�'!�'!�K?6��vo���������TH@�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�K?6�'!�'!�i\S�����vjb�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�SE;�'!�'!�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�ZK@�'!�'!�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�aQE�'!�'!�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�hWJ�'!�'!�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�o]O�'!�p6��r2��r2��r2��r2��r2��r2��r2��r2��r2��r2��r2��r2��r2��r2�p6�p6��v��v��v��v��v��v��v��v��v��v��v��v��v��v�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�p6�                                                                ��                                                          ��  OldCreateOrder	OnShowFormShow
DesignSize'� PixelsPerInch`
TextHeight TBevelBevel1Left Top Width'HeightNAlignalTopShapebsBottomLine  TLabelLabel1Left3TopWidthNHeightCaptionAnge &kommando:FocusControlCommandEdit  TLabelLabel2Left3Top8WidthWHeightCaptionAktuell katalog:  TLabelLabel4Left3Top"Width�HeightAnchorsakLeftakTopakRight AutoSizeCaptionP   Varning: Kör inga kommandon som kräver användardata eller dataöverföringar.  
TPathLabelDirectoryLabelLeft� Top8Width+HeightIndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TImageImageLeftTopWidth Height AutoSize	Picture.Data
�  	TPngImage�PNG

   IHDR           szz�   	pHYs  �  ��o�d  dIDATx�cd`�8� �cVpH)���_NMP�9�wG]m/��a :��:�:`��&T����g6M@u��U8]p��J�D�=������7/3���� E���6tu��#;�ܿ�p���]p��T�:���N@u���-]p��aTh�[��7.Gu���)]p��iT(k��w��Gu��*�(�Jb01�c�>w	��gh��/�:@VI,QW����� f��w����?Q���]Gu���X�	(�Ð���������W�	Sf3lݹ��x���$d�PHIJ0Tg3X���'Ϝgh������8�œ{���ê��ӕ�����������w�~Tq���P $*��HEY�����AOG�ߴu'CmS'U���3T��%YYYҒb����W�^�"�����b9|x�
���B`	-���U%���1�Y���g�T�/_�R�r�����x������6��jZΜ�@U�a�ۗO�`��K��3h��1�X�����_4�~~��� VVv�Y�����LL�tu��Q�H���o�;@D]���+=m����ۛ�7?���@ iC0�o    IEND�B`�  TMemo
OutputMemoLeft TopNWidth'Height;TabStopAlignalClientColor	clBtnFace	PopupMenu	PopupMenuReadOnly	
ScrollBarsssBothTabOrderWantReturnsOnContextPopupOutputMemoContextPopup  TButton	CancelBtnLeft�TopWidthKHeightAnchorsakTopakRight Cancel	Caption   StängModalResultTabOrder  THistoryComboBoxCommandEditLeft� Top	Width� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeCommandEditChange  TButtonExecuteButtonLeft�TopWidthKHeightAnchorsakTopakRight Caption   K&örDefault	TabOrderOnClickExecuteButtonClick  TButton
HelpButtonLeft�Top*WidthKHeightAnchorsakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick  TPngImageListImages	PngImages
BackgroundclWindowName&Copy log entries-console window outputPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?Cf���X�1&���Ӳþ`��e=��(�g���?���K��t���VC��w��?�,����(
>}��p��+���/�a`f�U����k�Ϫf(�u .�o��������W�+�_1��u�����������_�D��m؃-L�$���?�*��t�A����>2`�#�2�ه�I�+�Ϫg��₪i���Ʌs̬�3�}ހHhZ�vu$C�\�>��0�<g�\����Wg���oX�vMû���k�md@8���kO��;�1 �l@\����j���K~x��9LЁ��æ�g�V�A��]4 ������c@t�����i��F@������Y�����GZ3���fXP1���EA\��0�jH�*������]�&�(̊��o%â�X�D�,@	l��9Ò�x�DU���@Xښ� Ld8��h��    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
i  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?%�d@D�l�LYљ�7`ak
I�����%C���������́!�P3Հy�.�z°x�1�7�?��|<�����z�p5I�h�mJ����7Cq�
���2ؙh0�����ȹ[l�,��bX������0�b��_�n�����Ƞ�&����?���k�~���W�Nj=��������ÉKwn���%��o?��]��\`vZ�3�!|����y��o� �W�c�T�b�y���%d4�0�.,q��u�U�O0��3D�X�Ū&�b���+Cgq$܀����L��p��=��2�
�1��2\�������`���`1a>0;�̀�5	`���x��b7��  +!� "��p���hkU�xn�T&A �(��������e���8*��X�j���X�0��ߊf E��  O	��NV    IEND�B`� 
BackgroundclWindowName"Auto adjust size of console windowPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  2IDATx�c���?�y�u��mF���JI�=���n��M��:�b����O���/�g�+�*w��v���N
�,�g�Dfa�_<�a�����εs04����?�0@M�,�w�bg�X�"|�[WN#PT�c8�cX��#�$�·�����n`8��9 �>�w�<P� 	iE�Ӈ��%Lm1C��Լxza���4X���p��o_=E�'(�⼫g�`8Y�5�>��0���C��˧�lu]S�o_?#`ecg��ݸȠ���U����p>�<��/`( �h����`    IEND�B`�  Left�Top� Bitmap
      
TPopupMenu	PopupMenuImagesImagesLeft�Top�  	TMenuItemCopyItemActionEditCopy  	TMenuItemSelectAllItemActionEditSelectAll  	TMenuItemN1Caption-  	TMenuItemAdjustWindowItemActionAdjustWindow   TActionList
ActionListImagesImages	OnExecuteActionListExecuteOnUpdateActionListUpdateLeft�Top�  	TEditCopyEditCopyCaptionK&opiera
ImageIndex ShortCutC@  TEditSelectAllEditSelectAllCaption&Markera allt
ImageIndexShortCutA@  TActionAdjustWindowCaption   Anpassa &Fönster
ImageIndexShortCutJ@    TPF0TCopyDialog
CopyDialogLeftkTop� HelpType	htKeywordHelpKeywordui_copyBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption
CopyDialogClientHeight� ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize��  PixelsPerInch`
TextHeight TImage	MoveImageLeftTopWidth Height AutoSize	Picture.Data
�  	TPngImage�PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx���}Pe���!h�x�H$�^F���(��diYM�L��ț��d59���L6�$b�H�&h(�D`:9�"� ��	��������qw�t�77���>����=ϳ{��j��<(PUU;^E=EqK�j�ޛ�Bn;@���q�:vtt�������b���`0B�����;^!�7�e-B�^�(�5�����,�<vRN��B�yЎhi�s�����"\ B@9���/x�wB��hJH����L�i4������<_�G#��`6���3���� �a���$;�n'��g,֥y�w� >~!��<ڀ���s��~��rA�Htz�--T@ p��h�?�ѯc�gs��`2�d�*�$XN���=�q��I���4u�`Ѣ0�
ɀ9%���45�ǦCU�ݑ�ƀ΄n�QD<�ۯ���Mj|�3`TX��g���ӄ�?@0G<�A�����0�*���8}Z�ڛH�yv@\\�0!X���_�㪩���{���e?"J����c��%Л9|y����)�q�K�Z�4F�"��bPv@l�|q
�G��,W���e��{X���E8|�{?N������x�Ϙ��߭Ey�+o
1F��F�}����|�oA��y�`݈�)dDd��1Y��h΁��C��v��*�U�A��`�'���_�עQ[#&��˖\aki�2���8�T��'TbЇ�$���i�k��+�$�E�2�}��X��eq
�ƀ2`ʌ�d4�3���9M��6��*A���h����Y!��l@��HM۬����@L�K"��Q�KW�w�S�������da���c��$L
Q`V���55uh��d�����/V: �	�Z�ÈI���9u� �϶�}]��X�B�!�o�5XBr�xk�b�9�7�K��S�ajC��L(gOF�L���4�Z�QSTYvuk;%+�y��x������a9s�/Ցѡ�3��;U�"���Xl=�6�C��Z�0��s�AO�I�L>;��)$+��S(��4`$"z�*08$x��m���rj�>��o�J`o1�n�@ *G�[����F��G�ڷ��zP���4*�tHV`�"n_-N���y,��EO�>�8f��x��� ���x�� G��a��izD\oR'J�P�a�d��:��r����箟�yN�J��Î�:��� 
q"7�s"v\%͋��FOZ��.]ֵv��<��}�B��    IEND�B`�  TLabelDirectoryLabelLeft.TopWidth� HeightCaption)Copy 2 selected files to remote directory  TImage	CopyImageLeftTopWidth Height AutoSize	Picture.Data
�  	TPngImage�PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATx�ŕiPSW��{C�V��Ŵ��L�W�#�U��:ZG�-(���8���u�u	!@�mA� 00T��b���Tp�U! K"	f9��WÖ�eƓ�snN�����|_(B^f� ��5���Uk��)@9q���X�\Xc�a~�/w�Gc�5���� ��:#j�~�.��5��b�Fg@Ã�{T��:�B𱨀�1l�]&ǣ���;���E��[�B{O�h��)���Bb�����@�=�[����w@t��p�V���	`����l�e�{��-.:��m=��܃��~�x���_Χ��9����jzU:��u�{�y��� mK�� 6�(#i1�i�U��&�F�i��l1D/!����b �i�sk1u���h1I�A�R���
ޠ�1u�y��n_��u��c����Έ~bHY#@��B��c�(+�h��&�n�������'ҝ�B��Y��k_��Λ8�_�Y����W1u��1�X�M��Z�B�$�Ev�Z�SP�5���U���ǻ$�����&�n01( ,)�Hw�B�Bcܹ�*�}����̎�u��i e�y���T����6&AL�&�ED�g5��Q���,���ř�b��ē��x�6��F�*҉���P�x�v�YG��J�3ʹI�B`M��D�m�$V�Ǎ��Yq��p���i(��96��$�n�El�ǊG?;����m��"NV��m��g{N�8�953upp�gvC`z�XO��jH�!��O���Cd�>����ÂWN�w rۋee�ؾ�X�+�H�a���݈�a7pvw"n�4�w1��v6�0�S�ޯ�s�T֢.�1��Rd�X��ܙE��k�,�.�b'a/���4�A ��}�l�N���A�9��W0��6+�����Ӌ��{� ���*An;fb��\��p���HG�QUy5j7��:/�	��]�P��Qa��l�_/7w�)C� � V\�D ��N�
yP���+-�x�-��ӧ�"&ş�]*-GMD�	i�8���`0��l�����iq�ː�%�J�_�K9����!�s� ��]�zB]�9�O���eLǑ�A����Z��ׁ��s����B\Ċ-�oHт��@�j6�ލ�8��38s`�e��B��4=ȁ�E*���ÚyH:�������M��=[��7�E"_� &�,�0e�� � �P�e|��`�wx�j�Zo���h�\#��l��^��J�    IEND�B`�  TImageCopyUploadImageLeftTopWidth Height AutoSize	Picture.Data
/  	TPngImage�PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  |IDATx����Ow����bt:DZ"c$��mɲ� 4��͇=h�4�q�6�I�C%c@pBKA��fb��'�l��ln��x�'���B�~ww��X��?�\�z��}^����+E��Y�(J֠c�2���v�lQ�EY�{�޾
c"!e��W�Ң�wx�3Ni��� F�������8f�z��Л'݈_)�-��QF��e?���(�N�����ؼ��06>	���#F8D��=��7�D}$��I�'�a�vJ:~�`!,���k��=�+>J���qo�:5����^�=sd3�tfܼ7 �����!��sP>��m!���29#y���3h�������.@Jy��\�m6�$m��� ��M���o�j�Ɨ���Ҥm@N��7�4y;FY����i���vO��\��C��&+���Vy3��_gi�Qv|�'@j��
k�>�F��3�Uֈ��w\ ��"'��W�J}��he5Ή}�_g��P������.+��_UC������.�Ņ��� ��m�r��=�'��0�द���c�Eyy�������*+�	���N�����p��n�U�x1,4����B��cL��g�9Wjj���. ����ɵe�u�>�[V;C�~��(�������uB�%�3�Cg����%��"(L�jm� �����ɵ�d�:� 8��2�����C�"T�L�։ 1�5DN���T�4� ���OgEj�����R2�xqD}}� 8�WM���l2�$���G�4�(B�!X�6������*"'�)y��'?t���K�b�B)4��hj�^&�\˩蝛�p�6C"�F	j�ѓ-͍���Kĝk9�ϰ�%�X��@`P���Rz�Ǵǅ���$ �?���s-�&���,�"l#W+f? ������=��"�mu#ڮ5����d~��T�Nu�e^X,\\�F=�\�e$�G�q'an��m"��ߐ�r�u`���o��;#�a<���7���ō	�nu#�k{����b��V̌��B�� FM:<|���]<L;�,�u�AZ��k��S�  ��}�	���\������c�du��],[�e�Wb�Q���c}�g4�^�]�?�L����^��n���}�ʐ    IEND�B`�  TImageCopyDownloadImageLeftTopWidth Height AutoSize	Picture.Data
�  	TPngImage�PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx���{LSW��- ꘏��tnQ3�͹G�?���x+*��M����2�92�Z
��6�mq�F�`>��Ƕ8�RA)��*��E[�g���B�jz���4��9��>�w��\����(;��(A7핵
TSXl$R�f|b����&y���\������ihƻD������?o��!���t(�1�3;S ��3Æ��S�9��8�����[�=f�u�BcG�R�Q�5vĔ 9�_I�k1:�x5��P?��Лq�]�^����SdW�Bʲ"`��ȯ��ر_�X��A.���du^�S?@��HjJ�]eM�dv�f��{6�J�g1z�w�u9*r�y���6Au�0J�C�=@PP�"8=F����wH��N ���;Ԏ"1tf��8Z��	�}q� �u�TЩ�WrG2��^,����������~����Y�~�2 �jD́x`?X�S��n*a1�͋�(s�JΡ6?��^�v]�U�Ŭ�8�[#���mX��#��'�Ca�Y�l�9�-O��Mz��x��us��`я�����*����/L���7O�����?W׹�a.cZ9r7�o��fr�F�������o�Rx@V�ER�;�Q����b-��9>8u�g�`6Nd�D���R<��?�Y0���q"���j���v��@*����i�Na��a`�e/��h�s�M	x����.{p��;�4li� �;G$��0b�����k@�x*��WC���@�	�X�AÂ��X��<�}! �����~ͨ6���dm �܍6
��jɋ��&U��`�φ��\��As�`�kp{�S��bLd�߆;J���9@���k@�k�B���@�=��������[�Dp-�22)mX�N��1�	ӏ�D��6��@p�B�G�uY�r���k����c�!�� �x4���@�y@m���׀KT&�b#n2��2�0�tw��ge�2O��:M��0d��КE�]�������y[��	����4?�W5xh����|��#b�o��;�
Ni�6�e ��%�o��!��z�{qW~O)��{��J����T���H�pyf67%L*5Ϗ��[��G 8@R^-��
�����5~�#���
q����!�4�
�bN-FrB�3��\3���������V�mE�� E~�n=[��B�m75�d�i�� � ���Z�    IEND�B`�  TImageMoveDownloadImageLeftTopWidth Height AutoSize	Picture.Data
�  	TPngImage�PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx���{LSW�o�E|e:ԩ�
�%[�?f�"�"���|�#E`�L�.l�&��J�h6��Ő���:�g_��
}�׽���ֶt�p�X�!�7�������#"��U6� �M�x�@���5neQ�F�P(�A��c}�wt����GTĨ E��p�`0���Q�x�<�F#>|􄢤���G�z�hnV;v��$��b���D�S��-�!F�-ȧ�d20D�*�"����Fp�����;6iAb���?^C^^�ht �[м0@uM���s+r�4g9�EKK����������p���d��(���hh������D�$�U�k� 4ï����bs����RH��_���s��k�#^�@�3�8���~�.OBl�DPjj~
�T�#'���e��½a'۱�6'L���E�4�\81�1#�;���
ح�KN}��A�K�K��?au��y/�3ޏ:���;og#iڻ8���T,Em���\=9]�
��Ɓ���?���a ��au��a��
����:����!�E�z�(�C�J�D���!���!gv����v4���e��{������-8�����`3��y$3i�N�=���rG:
v��E�~'gw��� �Ҫzވ��RL�(��j\�Վ���#27G��SǱ`��g���ַ�mk�� ;O�J�}��A~�[�-:���͆��A�kN�g3W����92�M���_� ��>���� ������@���7�wx�xs _�]�n��9p&�N��e>9!�^�=$p��=��,ª� ���W��lV���ӱ$U�-ڥ킳���rbJ�L���Ƅ��&;�n؉���Aʿ�����7��فeiK������K�x-~�?2��p�Ȋ�GIa���N��6�d�
�����HO	��_���i���,�m�b��"L�L���5DY�&�C�y�
��:��&�̖�1��B�қُ}����)��9TM��7�hV�䪙X�qzX��3�eD�3MD� `��?偭���:ހ{�"��X�/;CGE�t�jj�<�Vz�(K��`V���@��uQ�N��V�GGK�n��|�Yb�El9p�(˲9��Mހcwaú�C�Z�נU����\r��+���/�BV榗~l{��k8DG�d�"g�r�S ���,l]�5��x�Ѩ�hU��'�-��Ek�p6�F�'��}�U�U���*��/.    IEND�B`�  TImageMoveUploadImageLeftTopWidth Height AutoSize	Picture.Data
?  	TPngImage�PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx����Ow���3� c$"�-Y���&qӹ�(N�a�����$��6����3J��4s����my�� ��zm��}{�У]��?쓴�\��}��s߻�˲�?�r(�5��H5u�f�-��&��\����8i�s�˷�hՌx `wk�O`b�Ư��y����� �~F��.��-ř���e?�g2�A������cߍ����Y1�D��%���q� ��[س�7c��t����~�a4㗎�2�s~�J�����Ŏ?�<��}�ѧ����g,����� sP~�kb��J��l<�Ar�F�1r�ͭ�9��?A�}��1%��bj�A^E�(�ɽ/�D[Q���(=�u����}�3r��eJ��a� ��<e�G��#l�Cg ?�c&����u #���)Qv�u� ��Aql&�; +�Gy�|��f�J��9pӦX8]y�[�@Y/*� �5�3_^��ܷ� ��*h���WCq|'�&���/��7��,����90v��WT����f��=� �V^�܁���\�X�<u�����q_H�X�&OGECB��|�H��2��m�=s�\�F�;� ����t.	(��ŉD�q�U��?���荂��4)h���I%yI����$��;x"$J�����t@��ZPT������~��ݡ�)��5^ f�YP����RY*w	ܫOgBNY"�6 <<b.�;����HMM��t���{I@��;(������?�lCXdB�"H(���B���y��{��@�Ƃ����.,|!���a %%�tw�
B��]��/ڰ&<!��A�-�hj����D���������a1X:�^�1�c��浦/ ҁ�����ǬȫB9��asg�^7���������H��z#���G�pV��6���dp���Z�0��pm���$q�,5�`�[.DK�"@R�n�<��8U;��J��u���q���T\x����1�ҺH�S����lv�V�C�H�bbL��.~��8��0���=@�\����n���x��WA����L��(u/b���C��\����n��?�����K�f�?r�l����*$�������M    IEND�B`�  THistoryComboBoxLocalDirectoryEditLeft.TopWidthtHeightAutoCompleteAnchorsakLeftakTopakRight TabOrder TextLocalDirectoryEditOnChangeControlChange  THistoryComboBoxRemoteDirectoryEditLeft.TopWidth�HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeControlChange  TButtonOkButtonLeftTop� WidthKHeightAnchorsakTopakRight CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeftWTop� WidthKHeightAnchorsakTopakRight Cancel	CaptionAvbrytModalResultTabOrder  TButtonLocalDirectoryBrowseButtonLeft�TopWidthKHeightCaption   &Bläddra...TabOrderOnClickLocalDirectoryBrowseButtonClick  	TCheckBoxQueueCheck2LeftToppWidth)HeightCaption1Transfer on background (add to transfer &queue) XTabOrderOnClickControlChange  	TCheckBoxQueueIndividuallyCheckLeft8ToppWidth� HeightCaption)   &Lägg till varje fil individuellt i könTabOrderOnClickControlChange  TButton
HelpButtonLeft�Top� WidthKHeightAnchorsakTopakRight Caption   &HjälpTabOrder	OnClickHelpButtonClick  	TCheckBoxNeverShowAgainCheckLeftTop� Width�HeightCaption$   &Visa inte den här dialogrutan igenTabOrder
OnClickNeverShowAgainCheckClick  TButtonTransferSettingsButtonLeftTop� Width� HeightCaption   Överförin&gsinställningar...TabOrderOnClickTransferSettingsButtonClickOnDropDownClick#TransferSettingsButtonDropDownClick  	TGroupBoxCopyParamGroupLeftTop5Width�Height2Caption   ÖverföringsinställningarTabOrderOnClickCopyParamGroupClickOnContextPopupCopyParamGroupContextPopup
DesignSize�2  TLabelCopyParamLabelLeftTopWidth�HeightAnchorsakLeftakTopakRightakBottom AutoSizeCaptionCopyParamLabelWordWrap	OnClickCopyParamGroupClick    TPF0TCopyParamCustomDialogCopyParamCustomDialogLeftvTop� HelpType	htKeywordHelpKeywordui_transfer_customBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption   ÖverföringsinställningarClientHeight�ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnCloseQueryFormCloseQuery
DesignSize�� PixelsPerInch`
TextHeight TButtonOkButtonLeft� Top�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  �TCopyParamsFrameCopyParamsFrameLeft Top Width�Height�HelpType	htKeywordTabOrder   TButton
HelpButtonLeftPTop�WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick    TPF0TCopyParamPresetDialogCopyParamPresetDialogLeftTopzHelpType	htKeywordHelpKeywordui_transfer_presetBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionCopyParamPresetDialogClientHeightClientWidth�Color	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize� PixelsPerInch`
TextHeight TLabelLabel1Left
TopWidthZHeightCaption   Förinställnings&beskrivningFocusControlDescriptionEdit  TButtonOkButtonLeft�Top�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft�Top�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TEditDescriptionEditLeft
TopWidth�Height	MaxLength� TabOrder OnChangeControlChange  �TCopyParamsFrameCopyParamsFrameLeftTop3Width�Height�HelpType	htKeywordTabOrder  	TGroupBox	RuleGroupLeft�Top[Width� Height�AnchorsakLeftakTopakRight Caption   Regler för automatiskt valTabOrder
DesignSize� �  TLabelLabel2LeftTopWidthOHeightCaption   Mask värdna&mnFocusControlHostNameEdit  TLabelLabel3LeftTopDWidthOHeightCaption   Mask an&vändarnamnFocusControlUserNameEdit  TLabelLabel4LeftToptWidthrHeightCaption   Mask &fjärrkatalogFocusControlRemoteDirectoryEdit  TLabelLabel5LeftTop� WidtheHeightCaptionMask &lokal katalogFocusControlLocalDirectoryEdit  TEditHostNameEditLeftTop$Width� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeControlChangeOnExitMaskEditExit  TEditUserNameEditLeftTopTWidth� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChangeOnExitMaskEditExit  TEditRemoteDirectoryEditLeftTop� Width� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChangeOnExitMaskEditExit  TEditLocalDirectoryEditLeftTop� Width� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChangeOnExitMaskEditExit  TButtonCurrentRuleButtonLeftTop� WidthIHeightCaptionAktuellTabOrderOnClickCurrentRuleButtonClick  TStaticTextRuleMaskHintTextLeft_Top� Width� Height	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaptionMasktipsTabOrderTabStop	   	TCheckBoxHasRuleCheckLeft�TopBWidth� HeightAnchorsakLeftakTopakRight Caption'   Välj automatiskt förinställning närTabOrderOnClickControlChange  TButton
HelpButtonLeftOTop�WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick    TPF0TCopyParamsFrameCopyParamsFrameLeft Top Width�Height�HelpType	htKeywordTabOrder  	TGroupBoxCommonPropertiesGroupLeft� Top� Width� HeightbCaption
EgenskaperTabOrder
DesignSize� b  TLabelSpeedLabel2LeftTopGWidthDHeightCaption&Hastighet (kB/s)FocusControl
SpeedCombo  	TCheckBoxPreserveTimeCheckLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption   Behåll tidsstä&mpelParentShowHintShowHint	TabOrder OnClickControlChange  	TCheckBoxCommonCalculateSizeCheckLeftTop.Width� HeightAnchorsakLeftakTopakRight Caption   B&eräkna total storlekParentShowHintShowHint	TabOrderOnClickControlChange  THistoryComboBox
SpeedComboLeftjTopCWidthUHeightAutoCompleteTabOrderText
SpeedComboOnExitSpeedComboExitItems.Strings	Unlimited10245122561286432168    	TGroupBoxLocalPropertiesGroupLeft� TopWidth� Height2Caption
EgenskaperTabOrder
DesignSize� 2  	TCheckBoxPreserveReadOnlyCheckLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption   Behåll skrivsky&ddParentShowHintShowHint	TabOrder    	TGroupBoxRemotePropertiesGroupLeftTop� Width� Height� Caption
EgenskaperTabOrder 	TCheckBoxPreserveRightsCheckLeftTopWidth� HeightCaption   Sätt fil&rättigheterParentShowHintShowHint	TabOrder OnClickControlChange  
TComboEdit
RightsEditLeft"Top*Width{Height
ButtonHint   Konfigurera filrättigheterClickKey@ParentShowHintShowHint	TabOrderText
RightsEditOnButtonClickRightsEditButtonClickOnExitRightsEditExitOnContextPopupRightsEditContextPopup  	TCheckBoxIgnorePermErrorsCheckLeftTopHWidth� HeightCaption   Ign&orera filrättighetsfelParentShowHintShowHint	TabOrderOnClickControlChange  	TCheckBoxClearArchiveCheckLeftTopbWidth� HeightCaptionRensa 'Arki&v' attributTabOrder  	TCheckBoxRemoveCtrlZAndBOMCheckLeftTop|Width� HeightCaption   Avlägsna BOM och &EOF teckenTabOrderOnClickControlChange   	TGroupBoxChangeCaseGroupLeftTopWidth� Height� Caption   Ändra filnamnTabOrder
DesignSize� �   TRadioButtonCCLowerCaseShortButtonLeftTop`Width}HeightAnchorsakLeftakTopakRight CaptionGemener &8.3TabOrder  TRadioButtonCCNoChangeButtonLeftTopWidth}HeightAnchorsakLeftakTopakRight Caption   I&ngen förändringTabOrder   TRadioButtonCCUpperCaseButtonLeftTop.Width}HeightAnchorsakLeftakTopakRight Caption	&VersalerTabOrder  TRadioButtonCCLowerCaseButtonLeftTopGWidth}HeightAnchorsakLeftakTopakRight Caption&GemenerTabOrder  	TCheckBoxReplaceInvalidCharsCheckLeftTopzWidth}HeightCaption   Ersätt '\:*?' ...TabOrderOnClickControlChange   	TGroupBoxTransferModeGroupLeftTopWidth� Height� Caption   ÖverföringslägeTabOrder 
DesignSize� �   TLabelAsciiFileMaskLabelLeftTopdWidth� HeightAnchorsakLeftakTopakRight Caption'   Överför följande &filer i textläge:FocusControlAsciiFileMaskCombo  TRadioButtonTMTextButtonLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption&Text (text, html, skript, ...)TabOrder OnClickControlChange  TRadioButtonTMBinaryButtonLeftTop/Width� HeightAnchorsakLeftakTopakRight Caption   &Binärt (arkiv, doc, ...)TabOrderOnClickControlChange  TRadioButtonTMAutomaticButtonLeftTopIWidth� HeightAnchorsakLeftakTopakRight Caption&AutomatisktTabOrderOnClickControlChange  THistoryComboBoxAsciiFileMaskComboLeftToptWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextAsciiFileMaskComboOnExitValidateMaskComboExit   	TGroupBox
OtherGroupLeftTopBWidth�HeightfCaption   ÖvrigtTabOrder
DesignSize�f  TLabelIncludeFileMaskLabelLeftTopWidth/HeightCaptionFilmas&kFocusControlIncludeFileMaskCombo  THistoryComboBoxIncludeFileMaskComboLeftTop$Width&HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder TextIncludeFileMaskComboOnExitValidateMaskComboExit  TButtonIncludeFileMaskButtonLeft;Top!WidthPHeightCaption&Redigera...TabOrderOnClickIncludeFileMaskButtonClick  	TCheckBoxNewerOnlyCheckLeftTopHWidth%HeightCaption!Endast &nya och uppdaterade filerParentShowHintShowHint	TabOrderOnClickControlChange  TStaticTextIncludeFileMaskHintTextLeft� Top:WidthiHeight	AlignmenttaRightJustifyAutoSizeCaptionmasktipsTabOrderTabStop	     TPF0TCreateDirectoryDialogCreateDirectoryDialogLeft�Top� HelpType	htKeywordHelpKeywordui_create_directoryBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSkapa katalogClientHeight� ClientWidthQColor	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSizeQ�  PixelsPerInch`
TextHeight TLabel	EditLabelLeftTopWidthUHeightCaptionNytt &katalognamn:  TEditDirectoryEditLeftTopWidthAHeightAnchorsakLeftakTopakRight 	MaxLength�TabOrder TextDirectoryEditOnChangeDirectoryEditChange  TPanel	MorePanelLeft Top2WidthQHeight� AnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneTabOrder
DesignSizeQ�   	TGroupBoxAttributesGroupLeftTopWidthBHeight� AnchorsakLeftakTopakRightakBottom Caption
EgenskaperTabOrder  �TRightsExtFrameRightsFrameLeftTop$Width� HeightWTabOrder �	TCheckBoxDirectoriesXCheckVisible   	TCheckBoxSetRightsCheckLeftTopWidth� HeightCaption   Sätt fil&rättigheterParentShowHintShowHint	TabOrder OnClickControlChange  	TCheckBoxSaveSettingsCheckLeftTop� Width-HeightCaption*   Använd &samma inställningar nästa gångTabOrder    TButtonOKBtnLeft[Top� WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft� Top� WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeft� Top� WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick     TPF0TCustomCommandDialogCustomCommandDialogLeft�Top� HelpType	htKeywordHelpKeywordui_customcommandBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionCustomCommandDialogClientHeightClientWidth�Color	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize� PixelsPerInch`
TextHeight 	TGroupBoxGroupLeftTopWidth|Height� AnchorsakLeftakTopakRightakBottom TabOrder 
DesignSize|�   TLabelDescriptionLabelLeftTopWidth9HeightAnchorsakLeftakTopakRight Caption&BeskrivningFocusControlDescriptionEdit  TLabelLabel1LeftTop@WidthXHeightAnchorsakLeftakTopakRight Caption&Eget kommando:FocusControlCommandEdit  TLabelShortCutLabelLeftTop� Width]HeightCaptionKor&tkommando:FocusControlShortCutCombo  TEditDescriptionEditLeftTop WidthfHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeControlChange  THistoryComboBoxCommandEditLeftTopPWidthfHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChange	OnGetDataCommandEditGetData	OnSetDataCommandEditSetData  	TCheckBoxApplyToDirectoriesCheckLeftTop� Width� HeightCaption   &Tillämpa på katalogerTabOrderOnClickControlChange  	TCheckBoxRecursiveCheckLeft� Top� Width� HeightCaption   Kör &rekursivtTabOrderOnClickControlChange  TRadioButtonLocalCommandButtonLeft� TopzWidth� HeightCaption&Lokalt kommandoTabOrderOnClickControlChange  TRadioButtonRemoteCommandButtonLeftTopzWidth� HeightCaption   &FjärrkommandoTabOrderOnClickControlChange  	TCheckBoxShowResultsCheckLeftTop� Width� HeightCaption!   &Visa resultat i terminalfönsterTabOrderOnClickControlChange  	TCheckBoxCopyResultsCheckLeft� Top� Width� HeightCaption&Kopiera resultat till urklippTabOrderOnClickControlChange  TStaticTextHintTextLeft"TopgWidthOHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	   &mönsterTabOrderTabStop	  	TComboBoxShortCutComboLeft� Top� Width� HeightTabOrder	   TButtonOkButtonLeft� Top� WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top� WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeft8Top� WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick   TPF0TCustomDialogCustomDialogLeft�Top� BorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSave session as siteXClientHeight)ClientWidthFColor	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenter
DesignSizeF) PixelsPerInch`
TextHeight TButtonOKButtonLeftETop	WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top	WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder   TButton
HelpButtonLeft� Top	WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick     TPF0TCustomScpExplorerFormCustomScpExplorerFormLeft� Top� CaptionCustomScpExplorerFormClientHeight�ClientWidthlColor	clBtnFace
ParentFont	
KeyPreview	OldCreateOrder
OnActivateFormActivateOnClose	FormCloseOnCloseQueryFormCloseQueryOnConstrainedResizeFormConstrainedResizeOnShowFormShowPixelsPerInch`
TextHeight 	TSplitterQueueSplitterLeft Top!WidthlHeightCursorcrSizeNSHintR   Dra för att ändra storlek på kölistan. Dubbelklicka för att dölja kölistan.AlignalBottomAutoSnapMinSizeFResizeStylersUpdateOnCanResizeQueueSplitterCanResize  TTBXDockTopDockLeft Top WidthlHeight	FixAlign	  TPanelRemotePanelLeft TopWidthlHeightAlignalClient
BevelOuterbvNoneColorclWindowParentBackgroundTabOrder  	TSplitterRemotePanelSplitterLeft� Top Height� CursorcrSizeWEAutoSnapColor	clBtnFaceMinSizeFParentColorResizeStylersUpdate  TTBXStatusBarRemoteStatusBarLeft Top� WidthlHeightPanels ParentShowHintShowHint	UseSystemFontOnClickRemoteStatusBarClick  TUnixDirViewRemoteDirViewLeft� Top Width�Height� AlignalClientDoubleBuffered	FullDrag	HideSelectionParentDoubleBuffered	PopupMenu&NonVisualDataModule.RemoteDirViewPopupTabOrder	ViewStylevsReportOnColumnRightClickDirViewColumnRightClick	OnEditingDirViewEditingOnEnterRemoteDirViewEnter
NortonLikenlOffUnixColProperties.ExtWidthUnixColProperties.TypeVisibleOnDDDragFileNameRemoteFileControlDDDragFileNameOnGetSelectFilterRemoteDirViewGetSelectFilterOnSelectItemDirViewSelectItemOnLoadedDirViewLoaded
OnExecFileDirViewExecFileOnMatchMaskDirViewMatchMaskOnGetOverlayDirViewGetOverlayOnDDDragEnterFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDQueryContinueDrag$RemoteFileControlDDQueryContinueDragOnDDGiveFeedbackRemoteFileControlDDGiveFeedbackOnDDChooseEffectRemoteFileContolDDChooseEffectOnDDDragDetectRemoteFileControlDDDragDetectOnDDEndRemoteFileControlDDEndOnDDCreateDragFileList%RemoteFileControlDDCreateDragFileListOnDDFileOperation RemoteFileControlDDFileOperationOnDDCreateDataObject#RemoteFileControlDDCreateDataObjectOnContextPopupRemoteDirViewContextPopupOnHistoryChangeDirViewHistoryChangeOnDisplayPropertiesRemoteDirViewDisplayPropertiesOnReadRemoteDirViewRead  TUnixDriveViewRemoteDriveViewLeft Top Width� Height� DirViewRemoteDirViewOnDDDragFileNameRemoteFileControlDDDragFileNameOnDDEndRemoteFileControlDDEndUseSystemContextMenuOnDDDragEnterFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDQueryContinueDrag$RemoteFileControlDDQueryContinueDragOnDDChooseEffectRemoteFileContolDDChooseEffectOnDDGiveFeedbackRemoteFileControlDDGiveFeedbackOnDDDragDetectRemoteFileControlDDDragDetectOnDDFileOperation RemoteFileControlDDFileOperationOnDDCreateDragFileList%RemoteFileControlDDCreateDragFileListOnDDCreateDataObject#RemoteFileControlDDCreateDataObjectAlignalLeftDoubleBuffered	HideSelectionIndentParentColorParentDoubleBufferedReadOnly	TabOrderOnEnterRemoteDriveViewEnter   TPanel
QueuePanelLeft Top$WidthlHeight� AlignalBottom
BevelOuterbvNoneTabOrder 
TPathLabel
QueueLabelLeft Top WidthlHeightIndentVerticalAutoSizeVertical	AutoSizeTransparent  	TListView
QueueView3Left Top-WidthlHeight_AlignalClientColumnsCaption	OperationWidthF Caption   KällaWidth�  Caption   MålWidth�  	AlignmenttaRightJustifyCaption
   ÖverförtWidthP 	AlignmenttaRightJustifyCaptionTidWidthP 	AlignmenttaRightJustifyCaption	HastighetWidthP 	AlignmenttaCenterCaption
UtvecklingWidthP  ColumnClickDoubleBuffered	DragModedmAutomaticReadOnly		RowSelect	ParentDoubleBuffered	PopupMenuNonVisualDataModule.QueuePopupSmallImagesGlyphsModule.QueueImagesStateImagesGlyphsModule.QueueImagesTabOrder 	ViewStylevsReportOnContextPopupQueueView3ContextPopup
OnDeletionQueueView3DeletionOnEnterQueueView3EnterOnExitQueueView3Exit
OnDragDropQueueView3DragDrop
OnDragOverQueueView3DragOverOnSelectItemQueueView3SelectItemOnStartDragQueueView3StartDrag  TTBXDock	QueueDockTagLeft TopWidthlHeight	AllowDrag TTBXToolbarQueueToolbarLeft Top CaptionQueueToolbarImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder  TTBXItemQueueEnableItemAction%NonVisualDataModule.QueueEnableAction  TTBXSeparatorItemTBXSeparatorItem203  TTBXItem
TBXItem201Action(NonVisualDataModule.QueueItemQueryAction  TTBXItem
TBXItem202Action(NonVisualDataModule.QueueItemErrorAction  TTBXItem
TBXItem203Action)NonVisualDataModule.QueueItemPromptAction  TTBXItem
TBXItem204Action*NonVisualDataModule.QueueItemExecuteAction  TTBXItem
TBXItem195Action(NonVisualDataModule.QueueItemPauseAction  TTBXItem
TBXItem194Action)NonVisualDataModule.QueueItemResumeAction  TTBXItem
TBXItem205Action)NonVisualDataModule.QueueItemDeleteAction  TTBXSeparatorItemTBXSeparatorItem201  TTBXItem
TBXItem206Action%NonVisualDataModule.QueueItemUpAction  TTBXItem
TBXItem207Action'NonVisualDataModule.QueueItemDownAction  TTBXSeparatorItemTBXSeparatorItem57  TTBXItem"QueueDeleteAllDoneQueueToolbarItemAction,NonVisualDataModule.QueueDeleteAllDoneAction  TTBXSeparatorItemTBXSeparatorItem202  TTBXSubmenuItemTBXSubmenuItem27Action-NonVisualDataModule.QueueCycleOnceEmptyActionDropdownCombo	 TTBXItem
TBXItem211Action,NonVisualDataModule.QueueIdleOnceEmptyAction	RadioItem	  TTBXItem
TBXItem225Action2NonVisualDataModule.QueueDisconnectOnceEmptyAction	RadioItem	  TTBXItem
TBXItem226Action0NonVisualDataModule.QueueShutDownOnceEmptyAction	RadioItem	   TTBXItem
TBXItem208Action*NonVisualDataModule.QueuePreferencesAction     TThemePageControlSessionsPageControlLeft Top	WidthlHeight
ActivePage	TabSheet1AlignalTopDoubleBuffered	ParentDoubleBufferedTabOrderTabStopOnChangeSessionsPageControlChange
OnDragDropSessionsPageControlDragDrop
OnDragOverSessionsPageControlDragOverOnMouseDownSessionsPageControlMouseDown 	TTabSheet	TabSheet1Caption	TabSheet1      TPF0TEditMaskDialogEditMaskDialogLeftqTopHelpType	htKeywordHelpKeywordui_editmaskBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionRedigera filmaskClientHeight�ClientWidth�Color	clBtnFace
ParentFont	
KeyPreview	OldCreateOrder	PositionpoOwnerFormCenterOnCloseQueryFormCloseQuery	OnKeyDownFormKeyDownOnShowFormShow
DesignSize�� PixelsPerInch`
TextHeight 	TGroupBox
FilesGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight Caption	FilmaskerTabOrder 
DesignSize��   TLabelLabel3LeftTopWidth=HeightCaption&Inkludera filer:  TLabelLabel1Left� TopWidth?HeightCaption&Exkludera filer:  TMemoIncludeFileMasksMemoLeftTop#Width� Height� AnchorsakLeftakTopakBottom Lines.StringsIncludeFileMasksMemo 
ScrollBars
ssVerticalTabOrder OnChangeControlChangeOnExitFileMasksMemoExit  TMemoExcludeFileMasksMemoLeft� Top#Width� Height� AnchorsakLeftakTopakBottom Lines.StringsExcludeFileMasksMemo 
ScrollBars
ssVerticalTabOrderOnChangeControlChangeOnExitFileMasksMemoExit  TStaticTextMaskHintTextLeft Top� WidthiHeight	AlignmenttaRightJustifyAutoSizeCaptionmasktipsTabOrderTabStop	   TButtonOKBtnLeft� Top�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeftTop�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeftVTop�WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TButtonClearButtonLeftYTop�WidthKHeightAnchorsakRightakBottom Caption&RensaTabOrderOnClickClearButtonClick  	TGroupBoxDirectoriesGroupLeftTop� Width�Height� AnchorsakLeftakTopakRight CaptionKatalogmaskerTabOrder
DesignSize��   TLabelLabel2LeftTopWidth\HeightCaptionI&nkludera kataloger:  TLabelLabel4Left� TopWidth^HeightCaptionE&xkludera kataloger:  TMemoIncludeDirectoryMasksMemoLeftTop#Width� HeighthAnchorsakLeftakTopakBottom Lines.StringsIncludeDirectoryMasksMemo 
ScrollBars
ssVerticalTabOrder OnChangeControlChangeOnExitDirectoryMasksMemoExit  TMemoExcludeDirectoryMasksMemoLeft� Top#Width� HeighthAnchorsakLeftakTopakBottom Lines.StringsExcludeDirectoryMasksMemo 
ScrollBars
ssVerticalTabOrderOnChangeControlChangeOnExitDirectoryMasksMemoExit   	TGroupBox	MaskGroupLeftTopqWidth�HeightLAnchorsakLeftakTopakRightakBottom CaptionMaskTabOrder
DesignSize�L  TMemoMaskMemoLeftTopWidth�Height4TabStopAnchorsakLeftakTopakRightakBottom 
BevelInnerbvNone
BevelOuterbvNoneBorderStylebsNoneLines.StringsMaskMemo 
ScrollBars
ssVerticalTabOrder       TPF0TEditorForm
EditorFormLeft;Top� HelpType	htKeywordHelpKeyword	ui_editorBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp Caption
EditorFormClientHeight}ClientWidthaColor	clBtnFace
ParentFont	
KeyPreview	OldCreateOrder
OnActivateFormActivateOnClose	FormCloseOnCloseQueryFormCloseQuery	OnKeyDownFormKeyDownOnShowFormShowPixelsPerInch`
TextHeight TTBXDockTopDockLeft Top WidthaHeight	AllowDrag TTBXToolbarToolBarLeft Top CaptionToolBarImagesEditorImagesParentShowHintShowHint	TabOrder  TTBXItemTBXItem2Action
SaveAction  TTBXItem	TBXItem16ActionReloadAction  TTBXSeparatorItemTBXSeparatorItem1  TTBXItemTBXItem3ActionEditCopy  TTBXItemTBXItem4ActionEditCut  TTBXItemTBXItem5Action	EditPaste  TTBXItemTBXItem6Action
EditDelete  TTBXItemTBXItem7ActionEditSelectAll  TTBXSeparatorItemTBXSeparatorItem2  TTBXItemTBXItem8ActionEditUndo  TTBXItem	TBXItem17ActionEditRedo  TTBXSeparatorItemTBXSeparatorItem3  TTBXItemTBXItem9Action
FindAction  TTBXItem	TBXItem10ActionReplaceAction  TTBXItem	TBXItem11ActionFindNextAction  TTBXItem	TBXItem12ActionGoToLineAction  TTBXSeparatorItemTBXSeparatorItem4  TTBXSubmenuItemEncodingCaptionKodningHint   Ändra filkodning TTBXItemDefaultEncodingActionDefaultEncodingAction	RadioItem	  TTBXItemUTF8EncodingActionUTF8EncodingAction	RadioItem	   TTBXItem	TBXItem13ActionPreferencesAction  TTBXSeparatorItemTBXSeparatorItem5  TTBXItem	TBXItem14Action
HelpAction    TTBXStatusBar	StatusBarLeft TopgWidthaPanelsCaptionLine: 2000/20000Size� Tag  Caption
Column: 20ViewPriorityPSize� Tag  CaptionCharacter: 132 (0x56)ViewPriorityZSize� Tag  CaptionEncoding: UTF-8 XViewPriorityZSize� Tag  ViewPriorityFStretchPrioritydTag   UseSystemFont  TActionListEditorActionsImagesEditorImages	OnExecuteEditorActionsExecuteOnUpdateEditorActionsUpdateLeft�Top8 TAction
SaveActionCaption&SparaHintSpara|Spara fil
ImageIndex ShortCutS@SecondaryShortCuts.StringsF2   TEditCutEditCutCaption	K&lipp utHint?Klipp ut|Klipper ut vald markering och flyttar det till urklipp
ImageIndexShortCutX@  	TEditCopyEditCopyCaption&KopieraHint,Kopiera|Kopierar vald markering till urklipp
ImageIndexShortCutC@  
TEditPaste	EditPasteCaptionKl&istra inHint0   Klistra in|Klistrar in innehållet från urklipp
ImageIndexShortCutV@SecondaryShortCuts.Strings	Shift+InsCtrl+Shift+Ins   TEditSelectAllEditSelectAllCaptionM&arkera alltHint%Markera allt|Markerar hela dokumentet
ImageIndexShortCutA@  	TEditUndoEditUndoCaption   &ÅngraHint%   Ångra|Ångrar den senaste ändringen
ImageIndexShortCutZ@  TActionEditRedoCaption   &Gör omHint&   Gör om|Gör om den senaste ändringen
ImageIndexShortCutY@  TEditDelete
EditDeleteCaption&RaderaHintRadera|Raderar vald markering
ImageIndex  TActionPreferencesActionCaption   &Inställningar...Hint:   Inställningar|Visa/ändra textredigerarens inställningar
ImageIndex  TAction
FindActionCaption   &Sök...Hint   Sök|Sök den valda texten
ImageIndexShortCutF@SecondaryShortCuts.StringsF7   TActionReplaceActionCaption   &Ersätt...Hint2   Ersätt|Ersätt den valda texten med en annan text
ImageIndex	ShortCutH@SecondaryShortCuts.StringsCtrl+F7   TActionFindNextActionCaption   Sök &nästaHint:   Sök nästa|Sök efter nästa uppkomst av den valda texten
ImageIndex
ShortCutrSecondaryShortCuts.StringsShift+F7   TActionGoToLineActionCaption   &Gå till radnummer...Hint/   Gå till radnummer|Gå till det valda radnumret
ImageIndexShortCutG@SecondaryShortCuts.StringsAlt+F8   TAction
HelpActionCaption   &HjälpHint   Hjälp editor
ImageIndex  TActionReloadActionCaption	La&dda omHintLadda om|Laddar om fil
ImageIndexShortCutR@SecondaryShortCuts.StringsF5   TActionDefaultEncodingActionCaptionAnsiXHint$Standard|Standard systemkodning (%s)  TActionUTF8EncodingActionCaptionUTF-8HintUTF-8|UTF-8 kodning   TPngImageListEditorImages	PngImages
BackgroundclWindowName	Save filePngImage.Data
k  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?%�d�B܆Ì6�hZ{��� [��q����2�����ܕ����a���/����/
���l�֭[�/
`����T��aB3^�V��;vlE5��Ӈ����!�(^1`��m��yx1���'��%k����{v��������_�� ����ph�NT�\<~(sgf�bĪ����];!^8zp���?~�%:Oރj���;��_�6��ѽ�Xۻ1|�	1`v<�7�/����~g���_~e���AD\��܉}�Xڹ2|��,�!G������<Kl Ƞ�5��$���O@5��ڙ������2�H�2tz~k���C��`1�r� � ��s�E�%�5�%�3���a�ehpz����nN����b p��!����L�w�g3H2H�_�ր�xG�F�L�  K��6B�    IEND�B`� 
BackgroundclWindowNameCutPngImage.Data

  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  aIDATxڝ�_HSQ����6�1_�BHP �T`0g0C�Az��-,�=&����X�z0T���H/i�� ��jnˠ@!	�nbX\��d�=�3MHY��p8�?����!8�l6G��F"���B �_|����yZ�R�J�p�(~�W�������/��&,������a|���(�{�A*
����N�r�"[Ų�����*��LLLΉ�i_���ȏ��5^����CZm�u�ǥ�8�~��,o��g�z��
 �E1@`�aѽ���7���ƞBWW'X,��b0<<�]Q��~��vtfw'"0���$��U�Os������,C(���3�����&������P��4�<Ǫ��j����_����c�mj:�y���4���Sgv��;r⓺�*�5�� mjһ��n�.��~6�
#��)��Z��5�/���SP*�K4}�-���GA�8�֭����\��-zD���V�k�J������Ul�P �)Kg�BGE�D��#B&!�mK3���w(�h+�fip6�����A�{rI�hE ���	���v��&�KDP(�~�~E�_q��x钱4�QVk�3|�O�O-���    IEND�B`� 
BackgroundclWindowNameCopyPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?Cf���X�1&���Ӳþ`��e=��(�g���?���K��t���VC��w��?�,����(
>}��p��+���/�a`f�U����k�Ϫf(�u .�o��������W�+�_1��u�����������_�D��m؃-L�$���?�*��t�A����>2`�#�2�ه�I�+�Ϫg��₪i���Ʌs̬�3�}ހHhZ�vu$C�\�>��0�<g�\����Wg���oX�vMû���k�md@8���kO��;�1 �l@\����j���K~x��9LЁ��æ�g�V�A��]4 ������c@t�����i��F@������Y�����GZ3���fXP1���EA\��0�jH�*������]�&�(̊��o%â�X�D�,@	l��9Ò�x�DU���@Xښ� Ld8��h��    IEND�B`� 
BackgroundclWindowNamePastePngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�cd@���]�����3L߸qm���	����?�#��]@Cmذ6�3��iǪ|��c�~0扌��-���79��Ǘ���cЛ��p���Ƿ�2 `�j�kx0�ۧ�Q$�}K���cL�ݧe�}��2�	�_f��3���.�(G.?dX���1&�_`C�8�1�ytŀ�ߓf�2|��E�ӗ�W�fX���9fVw�N!���_GQ��g2ì�`��Y�b��<��/�e�r�Ê]箂p�gxq�����a���/���;/�_{
f߹���n_AQ��_*��P�������æ�g ���2<�qE�2�4�Y�����j����m�`������E�Y�fWG2T����Hk����l��]>��`[&��(�w_�0���� H��3|z�Er�x9ì�h�����j.
�b��[����a�z��o��vAU�rF\�QU��3 
+�Ed��    IEND�B`� 
BackgroundclWindowNameUndo - internal editorPngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  cIDATxڝ��kRQǟs�L��9u��n�~̱�ʨ�6Al1�0X��z���{�Qob� �^hED4�
!iL�9�jfM�n���{o�J��.}�p~<���s��<��8���L+߇��ӰMoD���e�A�^T�������,J0T�ǡ	b2��pݡ;��`j� �/w����O_ �H�m��t��dǵ|b�eȭf�JK��ř� ��R�84�%�T�a�T���w�C�P����/�C�'�2沞 ,��j�ˬ� �SX7?�_0�7�Zh��{�(���\�������4D��0`K�y.��|�-B��}�")�� ��:��u����uQΦS���B�+��{h��I�RA�|� Z��HwR�U >�5v��c�\���n�m� �	Կd�佥P�ߔ+�	��Q�h�]�T["fA���0�/XIF>�Xv0:<�Y�75+�M�*ȥ�Bq�p-�������F�PK,����29���F���#*���\ :�OL,��b��S"�H�U*n@��f�cK�m��%R���&�Wb����$��e(�wǾ�2{5�тZ���u�G�ZF�J�Xih�����C��_���8�9�I4��    IEND�B`� 
BackgroundclWindowNameDelete - internal editorPngImage.Data
y  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڥ�KLQ�ϝ�N�@���R�����h1j���F�V���.\��n\��;I47�h(Y6PL�֐`+��R��t���̐"�������?�"B�O!	�gs�0�&^y����;�N�'{ �QBQ�����o�ļ���]	�t:��~�[|�k7P��ͧu:=�'���m �Y�Y�f��g>�LN8���N�zg4[��j���jdiD����ŝ��#@�l%A`���ø�dQ���Gs���d���y���SI�m�:ڛ�uuX�!խ��.�jj��hH&6 �����lY*k�R�"���0��i~ *��.�l�>R��Wmյ@3$6� CAQ	��Eaq!�9�0=>����.g��6˪�Y�A�`�^b3.���}��������H3��� �Rk�^<�"�^��� =�������a��[k(V�!���$P,��hx:�4���K�����P��Kkbd���ٟ%��ŮQkt]�	�U>մ�|}��ɹ*Y�S�h��l6#����Ѕ�#�5�*��"Ɋ�ɛ�1�yB�������JTj`������5/?�X�E>s̗-m�^������C�,N��]���c��a+�`���ݧ\��n'���2�P�Jx!.�w2�ov�ĕ��q>����g:v���0�qޞ�����Y����d���rb³)its����5    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
i  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?%�d@D�l�LYљ�7`ak
I�����%C���������́!�P3Հy�.�z°x�1�7�?��|<�����z�p5I�h�mJ����7Cq�
���2ؙh0�����ȹ[l�,��bX������0�b��_�n�����Ƞ�&����?���k�~���W�Nj=��������ÉKwn���%��o?��]��\`vZ�3�!|����y��o� �W�c�T�b�y���%d4�0�.,q��u�U�O0��3D�X�Ū&�b���+Cgq$܀����L��p��=��2�
�1��2\�������`���`1a>0;�̀�5	`���x��b7��  +!� "��p���hkU�xn�T&A �(��������e���8*��X�j���X�0��ߊf E��  O	��NV    IEND�B`� 
BackgroundclWindowNameDisplay preferences windowPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  JIDATx�u�{hYƿ;���S��M�*q׵�U�ڭ������u]�ڦ��c�e��������U�����J���
Q�'��R|���C-kk���mb��13��f�J������9����DY�s�
R��黦�[wp�:�1)�T+�R�C��5_���QQ�q½;gxXB����Wa��-Y�,9S���v`D y��7��~���-I��~W��Mu�j����}����X��h�d�B��{&b,�xj�4��r�/?̝�Z[�z�
��X:^cHa6����������q�D��O��A��&|����fQJ��ߎ�23L�䄖�TP�0x���A�0��&Ga�(�i?�o����i�T���D��E��TU���n4?~���q�k�*�Nd÷���_+W���̜�5���w��SX�/�l6��)�Aܼ�7����r��?K�ݻ(��.���s8T6&r�d�H���ǅ�	��<�d��$p��yQ8Z���|��EDQ��+8u�B$�ʓ���%ҹlI�`�	.�B�P�T��y�@��P�*{Η���%��U�=����<�c�r�M1Mϛ��)����Ez�o��S� �r,�s��� �,�s�F��Ȳ���݃z��O?ڨ�H`�ϋ̼� ��ǲ�e))zز-Z�o�}H1�p��dE�z��he��u�֬����F0��f�W'�^:M,�H7�CFz������@�%��򨫜�i����#����I%�?A�]����W=�T�:�`�p���$�Ƣ�>�0X�y�8%���Q���9i=�����ks����#����`E��VE�ț΍Z���Q��M?����䷆�u{ƪ{�/m�m$yL    IEND�B`� 
BackgroundclWindowNameFind text - internal editorPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  FIDATx�cd�55��@��=r��u[Br���g`DR���#�AQI�aѴN�"9~I%=}C��;���P�o��B]Ë��:��f�X��!M��r`���y~��w�W�i��.`@ۗN@�>�����Ν����s��m���l��p��M����1��Z�U��2��-f��� �0l�w����o�=�ze���f���f���'܀3���V��|j?Ã��'ܺu����Fv>*�&(.�cPW�f�dcax�����/���ܻq��ک��n޼fͨ����R��B�	����*l�̷�u�4Tn�}�p��i����޽{�H���嶒�)���4ý���\9�����;w����F�R��S=U���/3�;���ë��@����q�������Dy�1�H�0\�z����S��Y4 �<ЀhP<Tҳ�s��F'X��g.���������oܸ&Ϩ�o�����<�!�������3���/]8���P�_VQ��To�{����/}-%����uz�������݃˯���Rph��h:4��<� KFP��  ,/�A�x    IEND�B`� 
BackgroundclWindowNameReplace textPngImage.Data
i  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�cd�l���Y7����M`f"#�<0����#��'� l6�h� �P�\ 0`.����R��?w�ea�|� ������+�=��Ee�J�8���$cק=:��߻���z�����a��a9k��_���_�t�w66�{K.3������������}�b�˖���R���_��+��c@???;;ûw�ﱲ�JHH�s=��0����9P�[o���yRLT����������������s;�?�X���f��&222̃1$�CU>f�bi�aaav �`�|�گ��?	>���9f���O����3@��������"7;;;�����������Ar�B6 ���h�s]c���#�������{����uG�Nf���rQk����;��9��̰�������p�
b��^��� �%�����    IEND�B`� 
BackgroundclWindowName	Find nextPngImage.Data
P  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڍRyH�a�}N��Gba���v977�u�QxdA�E)�H�Z៕)�����A%�`�BA���i��y�sΉό��N�����ف?xy���=���}	,C 5�WȲ���O���H�B��!yxx��$+�u	�,MOk��U#�����)�O~E�m%J/���c��׊#�b��������+�����E��;��d��w~"��"]�=BbS,��]���?p��~s�ܟ��7*��hO�x�\�7��<:����V|�(ד�Ĭ
T�_��P~��,ХjĠ�C�N�9�t�H����XnՁ����'ض���"�z;Уz�B/3�
EE�\���a���Aؠ��:����Z ��r�<���+�_��z��j�ϙ�z}w?÷�4��i15kB�Y9>�_�RQ#U*]�|S؎Ί����#�Y���IH|ɛ����kj�e�ɉY��zH����E^�Ը�<))�=���e�WJlB:��nF{w?�rN�x�[�~b��r��ñ�7Ρ��=$�3/GL��4�;*:�~*�@YA�����`gk�-�|�>,�
��0�#�e����Y'�JZm���3.P;80_U;0�q2?��Ъ���%sCU��FF���,w�D8��O@�F�8�۝�.Q��nƇ�X'|��AaEP)��x�J��4&�����    IEND�B`� 
BackgroundclWindowNameGo to line numberPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  5IDATx�c���?%���ѻ�d�PH���F�?ï?ę�7a�i����,`(�u���D;��~�
���30����\��g��� �o?���	��700b�y�:� �7����-ˎ��g�PԿb����/��ܾ����S��pWc)��OX�0����������G�Neؼ'�f�/J��bwAi����$A���F>��[�}�W'��,�l@̺�@�@�`��i߬�h�w_��+Q�Al���j���"��(Ԋ�݀�@b�|!�U��Q���Gz^�87Rj  ���qx    IEND�B`� 
BackgroundclWindowNameOpen online documentationPngImage.Data
i  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�mSKLQ=3�ϔ��P@
���E���2��Ѱ�HPQ�G�l\�V?$�� @4ą���L�5�������Ng|�P�[����s�}��m��a��Pb�@�E���R�GA�^:^��m�S�^*��!V�H�Ȯf��Ӛt�JV�b\��+K�;5���@}4!�yx4]�U�k*��n�!��x�J�,��<5p�M"��|$"5�"�@Q��3��p�XX&e��&q�5MЪ�fx0`âXF&���A���l_���4X�@i-,�G�4�d�w\���\�_��ǣ�@P�1��A�pL|#;WA��gd�鳌RvK�m[��a�~�%d5��=]���.�M�Uz�Xq�w�ak�y�E�Tm�*i�̡t|����tϠ�V%,Ez\x���RL�E�0���(���x�����p��b��d���2����H*sLI;-��tX��#&���1�՟�������r�wY�
6E�EKX��nG
�F��0c�.Q��n��)�l��d��çb!�����T#-*��(��6�ͅA+Gs�\J�����
�H�s�]JV}Y��#��~ތ��]SIq��"��j����J�ʫ����M���d��*ebo/��ꘚ�&��Qɟ�íl��^���$L����#kA����ñ�I?��U�8����VJD�4m��D
�d��3�w��V�_l�'|=&.    IEND�B`� 
BackgroundclWindowNameReload filePngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  nIDATxڍ�]H�Q��6Ge6����,���E؅Q�2�ӥ�H7eN3�ۖ���.b4}3��o�&]ɊP�>�p�+A��s�6���A��P��꜇���s8�p!(��!X58ܵ�$ma�38�e���5/�㢳�x�w�5��o�z=2���0�J�s�+>ע��9]�|�����!��I���pY�Mt�,�}+Qkx��]���m�Ö:YJ�Uv�����g�E��_V��$��~	<�1��+!�$����R�.Ut����܇��F$=&��a{��.���[�����M�,���6r=�����gڶ͎��"��L�/r�4���@���з�1��]rv�[�?���B;�՝h��Y@B].��<T��I�,�C��`�ly���[V��X�£�%]�ֶ�"�2�� q73Eg�2Qt���WzK݊f��2ʞ���, �چ��-�ݸ��y����X��d��"�ĥ��� A-���#0O�<_�ߑ�-b�����#��M��t��R��%4��rq�D!�p�f�z�N��G|�.���N��O�:����Z��i�z����>�Y�S�
 m��p�V��?�.�w�    IEND�B`� 
BackgroundclWindowNameRedoPngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  [IDATx�c���?###6�ట���?�b*��D��`g����%�ψb@C��=��`6���s������L����3K�0�?����o�H�����+;�VAa;e~A���/_�<y�������hj��\�r���� Fb7l����PV�d���û�����3��3���3�}��P\RZ����]�(Į����ݢgd�����;7/�����F�(eu1q)x8�<�� ������x���^8�����&��]U��,����IEM	Aa1��N�G3 n�{M+���^3<}t{��Łq I���Kɫh�J����31��a`����]�����?X4	b���@�#~O�_�o�l�W%MS�o_0�}���ᒀ2 �)6�R�`ffex����?̺����!� ��Ŝ�<=�@�~����0����`i�	�\�����_�˼|B*\<?|c���=ÿ��n����)P��K�vc5 ���+���p���[���,����!���2�#�_�{��na5 ����gf������&ffPB˃\4��ޢ�=8���LL�@%6@y -T�Y�`,w�@	  �7�_�!W    IEND�B`�  LeftTop8Bitmap
      TTBXPopupMenuEditorPopupImagesEditorImagesLeft�Top�  TTBXItemUndo1ActionEditUndo  TTBXItem	TBXItem18ActionEditRedo  TTBXSeparatorItemN1  TTBXItemCut1ActionEditCut  TTBXItemCopy1ActionEditCopy  TTBXItemPaste1Action	EditPaste  TTBXItemDelete1Action
EditDelete  TTBXSeparatorItemN2  TTBXItem
SelectAll1ActionEditSelectAll  TTBXSeparatorItemN3  TTBXItemFind1Action
FindAction  TTBXItemReplace1ActionReplaceAction  TTBXItem	Findnext1ActionFindNextAction  TTBXItemGotolinenumber1ActionGoToLineAction  TTBXSeparatorItemTBXSeparatorItem6  TTBXItem	TBXItem15ActionPreferencesAction       TPF0TEditorPreferencesDialogEditorPreferencesDialogLeft/Top� HelpType	htKeywordHelpKeywordui_editor_preferencesBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionEditorPreferencesDialogClientHeightgClientWidth�Color	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize�g PixelsPerInch`
TextHeight 	TGroupBoxExternalEditorGroupLeftTop� Width�HeightIAnchorsakLeftakTopakRight CaptionC   Alternativ extern editor (påverkar bara redigering av fjärrfiler)TabOrder 	TCheckBoxExternalEditorTextCheckLeftTop-WidthQHeightCaptionH   Tvinga fram textöverföringsläge för filer redigerade i extern editorTabOrder  	TCheckBoxSDIExternalEditorCheckLeftTopWidthQHeightCaptionA   E&xtern editor öppnar varje fil i ett separat fönster (process)TabOrder    	TGroupBoxEditorGroup2LeftTopWidth�Height}AnchorsakLeftakTopakRight CaptionEditorTabOrder 
DesignSize�}  TRadioButtonEditorInternalButtonLeftTopWidth� HeightCaption&Intern editorTabOrder OnClickControlChange  TRadioButtonEditorExternalButtonLeftTop-Width� HeightCaption&Extern editorTabOrderOnClickControlChange  THistoryComboBoxExternalEditorEditLeft TopEWidthHeightAutoCompleteAnchorsakLeftakTopakRight TabOrderTextExternalEditorEditOnChangeControlChangeOnExitExternalEditorEditExit  TButtonExternalEditorBrowseButtonLeft1TopCWidthKHeightCaption   B&läddra...TabOrderOnClickExternalEditorBrowseButtonClick  TRadioButtonEditorOpenButtonLeftTopaWidth� HeightCaption&Associerad applikationTabOrderOnClickControlChange   	TGroupBox	MaskGroupLeftTop� Width�HeightIAnchorsakLeftakTopakRight CaptionAutomatiskt val av editorTabOrder
DesignSize�I  TLabel	MaskLabelLeftTopWidth� HeightCaption/   Använd den här editorn för &följande filer:FocusControlMaskEdit  THistoryComboBoxMaskEditLeftTop'WidthoHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder Text*.*OnExitMaskEditExit   TButtonOkButtonLeft� TopFWidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� TopFWidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeft?TopFWidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  	TCheckBoxRememberCheckLeftTop.WidthQHeightAnchorsakLeftakBottom Caption   &Kom ihåg den här editornTabOrder    TPF0TFileFindDialogFileFindDialogLeftoTop� HelpType	htKeywordHelpKeywordui_findBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp CaptionFindXClientHeight�ClientWidth2Color	clBtnFaceConstraints.MinHeight� Constraints.MinWidth�
ParentFont		Icon.Data
~           h     (                 @                                      saR�s`R�s`R�s`R�saR�    saR�s`R�s`R�s`R�saR�                    s`R�������������s`R�    s`R�������������s`R�                    50.�)&&�)&&�)&&�50.�    50-�)&&�)&&�)&&�50-�                    )&&�QD:���o�����)&&�    )&&縬����o�QD:�)&&�                    *''�MB;��xg���}�*''�    *''���}��xg�MB;�*''����������������"c��B:5�]PG�KFD�"_{����#]x�KFD�]PG�B:5�(%%Z�������������������Ow��)&&�)&&�)&&�)&&�)&&�)&&�)&&�)&&�)&&�)%%����:���7���7���7���.^m�eVL�������o����������ym���o�����eVL�)&&����V���I���I���H���>���E<7�������o�)&&�)&&�)&&���o�����E<7�+''T���e���N���N���N���K���.>B�)&&�)&&�)&&�+01�)&&�)&&�)&&�)&&�+++���s���T���S���S���S���R���)&&�����)&&�Q���)&&�����)&&�        ���������������������������UWW�)&&�SUV�����&;F�)&&�)&&�        ������������������������������������                ���4���4���4���4���4���4���4���4���4���4������                ���1���A���A���A���.���������������������                �������������������                                    �   �   �   �   �                                      �  
KeyPreview	OldCreateOrderPositionpoOwnerFormCenterOnCloseQueryFormCloseQuery	OnKeyDownFormKeyDownOnShowFormShow
DesignSize2� PixelsPerInch`
TextHeight 	TGroupBoxFilterGroupLeftTopWidth�HeightAnchorsakLeftakTopakRight CaptionFilterTabOrder 
DesignSize�  TLabel	MaskLabelLeft1TopWidth/HeightCaption	&Filmask:FocusControlMaskEdit  TLabelRemoteDirectoryLabelLeft1TopGWidth0HeightCaption   Sö&k i:FocusControlRemoteDirectoryEdit  TImageImageLeftTopWidth Height AutoSize	Picture.Data
�  	TPngImage�PNG

   IHDR           szz�   	pHYs  �  ��o�d  =IDATx�ŖL�eǿ������:���.�011��p!舻�\�T2��uS+Vkɼ�V8+A�i	z�@�wx!؄̚����x��8�`�����{����mϞ�}~���>����{'��l��Eáa���V<����z0M*=t�>% UE⏣�/�K��s
��|����j�N:�����3���M)���ن�p�q�n�'f��<� UE�1��\<��Wl�M���c���^�/ F�5f��iԉ6��	<�Y��YaS
p�Z�0���3^ YA�&�>\�`_�w���x��PW���cM~ ��% G�pˏ�q.���~ �ˁ�c���\�`I�W6���#7��? yG��3��~Z.-�����lWPptJ�5Bs��z��B�\�
d?��5���do�7��u<�AX^�Y��B�\V�:s�V�<������G�	�F0�#G^�{����=������Z|$�Q��+͆�@.���&����-�XI^�^�On� ��@ ������� KV�qGk�R�z���LzJ��XB��!�6t�wb�漨6��� -)��n�`��|߈��Qط}-�3��Z�R(/h`1Ѹ�<	�_77�0_� �����|��ÊO�Q�����n �rN}I�i���{���ZA�w;+�����٦rX��ai�� 22OH� ������.lް��u�͗�7�0I,��g�`������u�SJ*������q~�����f�ap�~�,sX���ry
�x�{sq)�HNx�߁��o4~WC�n���ph�G+��&wӨ/(10�?g$�(@/�f��x�v�E�t����:y����=&T��;W"z��W�ݩM�e�X�zX�<���u�����x�7]E7MCU_�?:Z�!��L�.*晌�򗑑�MW~��dk������@4�J�\/JM�Bl�"Gp��2RZT���n �q��>��c��원9s�Uw��Մ����=n�5[�bđ�;��7�HWۡ���X��5��łMjj
)�SX$y����Z�ؘ�j&�&S"������89�Dz`R�_ѹi?�X�    IEND�B`�  THistoryComboBoxRemoteDirectoryEditLeft1TopWWidth�HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeControlChange  THistoryComboBoxMaskEditLeft1Top$Width;HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder TextMaskEditOnChangeControlChangeOnExitMaskEditExit  TStaticTextMaskHintTextLeft� Top;WidthtHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	Mask&tipsTabOrderTabStop	  TButton
MaskButtonLeftrTop!WidthPHeightAnchorsakTopakRight Caption	&RedigeraTabOrderOnClickMaskButtonClick   TButtonCancelButtonLeft�Top+WidthPHeightAnchorsakTopakRight Cancel	Caption   StängModalResultTabOrder  TButtonStartStopButtonLeft�TopWidthPHeightAnchorsakTopakRight Caption&StartXDefault	TabOrderOnClickStartStopButtonClick  TButton
HelpButtonLeft�TopKWidthPHeightAnchorsakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick  TIEListViewFileViewLeftTop� Width�Height� AnchorsakLeftakTopakRightakBottom ColumnClickFullDrag	ReadOnly		RowSelect	TabOrder	ViewStylevsReport
OnDblClickFileViewDblClick
NortonLikenlOffColumnsCaptionNamnWidthP CaptionKatalogWidthx 	AlignmenttaRightJustifyCaptionStorlekWidthP Caption   ÄndradWidthZ  MultiSelectOnSelectItemFileViewSelectItem  
TStatusBar	StatusBarLeft Top�Width2HeightPanels ParentShowHintShowHint	SimplePanel	  TButtonFocusButtonLeft�Top� WidthPHeightAnchorsakTopakRight CaptionF&okusModalResultTabOrderOnClickFocusButtonClick  TButtonMinimizeButtonLeft�Top+WidthPHeightAnchorsakTopakRight Caption	&MinimeraTabOrderOnClickMinimizeButtonClick   TPF0TFileSystemInfoDialogFileSystemInfoDialogLeft@Top� HelpType	htKeywordHelpKeyword	ui_fsinfoBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption#Information om server och protokollClientHeight�ClientWidthsColor	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnShowFormShow
DesignSizes� PixelsPerInch`
TextHeight TButtonCloseButtonLeft� ToplWidthKHeightAnchorsakRightakBottom Cancel	Caption   StängDefault	ModalResultTabOrder  TButton
HelpButtonLeftToplWidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TPageControlPageControlLeft Top WidthsHeight`
ActivePageProtocolSheetAlignalTopAnchorsakLeftakTopakRightakBottom TabOrder OnChangePageControlChange 	TTabSheetProtocolSheetCaption	Protokoll
DesignSizekD  	TGroupBoxHostKeyGroupLeftTop� Width_Height)AnchorsakLeftakRightakBottom Caption$   Nyckelfingeravtryck till värdserverTabOrder
DesignSize_)  TEditHostKeyFingerprintEditLeft
TopWidthNHeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFaceReadOnly	TabOrder TextHostKeyFingerprintEdit   	TListView
ServerViewLeftTopWidth_Height� AnchorsakLeftakTopakRightakBottom ColumnsAutoSize	CaptionArtikel AutoSize	Caption   Värde  ColumnClickDoubleBuffered	MultiSelect	ReadOnly		RowSelect	ParentDoubleBuffered	PopupMenuListViewMenuTabOrder 	ViewStylevsReportOnContextPopupControlContextPopup  	TGroupBoxCertificateGroupLeftTop� Width_HeightHAnchorsakLeftakRightakBottom CaptionCertifikatets fingeravtryckTabOrder
DesignSize_H  TEditCertificateFingerprintEditLeft
TopWidthNHeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFaceReadOnly	TabOrder TextCertificateFingerprintEdit  TButtonCertificateViewButtonLeft
Top%WidthyHeightCaption   &Fullständigt certifikatTabOrderOnClickCertificateViewButtonClick    	TTabSheetCapabilitiesSheetCaption   Möjligheter
ImageIndex
DesignSizekD  	TGroupBox	InfoGroupLeftTop� Width_HeightrAnchorsakLeftakRightakBottom Caption   Övrig informationTabOrder
DesignSize_r  TMemoInfoMemoLeft	TopWidthMHeightWTabStopAnchorsakLeftakTopakRight 
BevelInnerbvNone
BevelOuterbvNoneBorderStylebsNoneColor	clBtnFaceLines.StringsInfoMemo 
ScrollBarsssBothTabOrder WordWrap   	TListViewProtocolViewLeftTopWidth_Height� AnchorsakLeftakTopakRightakBottom ColumnsAutoSize	CaptionArtikel AutoSize	Caption   Värde  ColumnClickDoubleBuffered	MultiSelect	ReadOnly		RowSelect	ParentDoubleBuffered	PopupMenuListViewMenuTabOrder 	ViewStylevsReportOnContextPopupControlContextPopup   	TTabSheetSpaceAvailableSheetCaption   Tillgängligt utrymme
ImageIndex
DesignSizekD  TLabelLabel1LeftTopWidthHeightCaption
   &Sökväg:FocusControlSpaceAvailablePathEdit  	TListViewSpaceAvailableViewLeftTop(Width_Height� AnchorsakLeftakTopakRightakBottom ColumnsAutoSize	CaptionArtikel AutoSize	Caption   Värde  ColumnClickDoubleBuffered	MultiSelect	ReadOnly		RowSelect	ParentDoubleBuffered	PopupMenuListViewMenuTabOrder	ViewStylevsReportOnContextPopupControlContextPopup  TEditSpaceAvailablePathEditLeft8Top	Width� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeControlChangeOnEnterSpaceAvailablePathEditEnterOnExitSpaceAvailablePathEditExit  TButtonSpaceAvailableButtonLeft TopWidthcHeightAnchorsakTopakRight CaptionKon&trolleraTabOrderOnClickSpaceAvailableButtonClick    TButtonClipboardButtonLeftToplWidthyHeightAnchorsakRightakBottom Caption&Kopiera till urklippTabOrderOnClickClipboardButtonClick  
TPopupMenuListViewMenuLeft� Topb 	TMenuItemCopyCaptionK&opieraOnClick	CopyClick    TPF0TFullSynchronizeDialogFullSynchronizeDialogLeftmTop� HelpType	htKeywordHelpKeywordui_synchronizeBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSynkroniseraClientHeight�ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize�� PixelsPerInch`
TextHeight 	TGroupBoxDirectoriesGroupLeftTopWidth�HeightwAnchorsakLeftakTopakRight Caption	KatalogerTabOrder 
DesignSize�w  TLabelLocalDirectoryLabelLeft1TopWidthJHeightCaptionL&okal katalog:FocusControlLocalDirectoryEdit  TLabelRemoteDirectoryLabelLeft1TopDWidthWHeightCaption   F&järrka&talog:FocusControlRemoteDirectoryEdit  TImageImageLeftTopWidth Height AutoSize	Picture.Data
�  	TPngImage�PNG

   IHDR           szz�   	pHYs  �  ��o�d  dIDATx�Ŗ{lSUǿ�]o[�G�l��Qb�и�(b�l1��m>�H܀�E2�-�4f	1�h�?�5D��R4��i���[�Y�u�n��֕�k{o{��-H��v�.�����������<n�ύ�q�fЩ�iB�Z/-%������0�_�syG
K���?$)�3�K����S����TiT%�>*cլ����h��'�?����[�_S
p�!�[���uw��M(���y��_ZM�x ��y}�~�d3�t��~���౲�
��y[b�u��� 嵿/�����I ^�
p�%����H��g<֞��g��9w%ђn��;� �|��͹�|u�FS���}b��D�Q��t)	��w�)	���Z)��9�9P�j�r���IR��Cs����s.(����پq\���� c��.¦�lh.��Z�g����@���h����%|�oEo �C&+�sB�4�ٙP+UP�Yp��S��O�b/.*����`�^��~�c'��<��U��YK2@8@�*��͢j�r%���v���y���� {wP�?�{�c�o�/V|7�	=���-���kҋe+�a�]��LS� �0��3'% ���K�7�����q���k�4�yآ���f�������Pt_Q�%�Q�X���? �gK�cS	�)8b��>S��9�Q�V/���Q�֮��7�b��T�D/ %��9^*$���Pz��kVC��2l�3r4~z<���<�O��$�bu׃"*�#�qK� ��ٛ0�X�����~���L+v@K��L;�ؔ� r�K��^�{��r"�x.t���r7������& �'�c<�����t��I��j�t�f�y
�?؇+W�� nz�a���NO������|J �ۺ+d�@�/�1<<� 0���ɑ�� �����ș�HX��p��q5% ;���/���z{za�Dhg��G��(t ��?�_�x&eS����B����7��������nIFIwƸ��[��7X�<)���e6O�e&�,Y��xi6X��&�����s̍ '�R�[�S��0Z�4�/�f�*
RF��K���^����-�u��R5�@*��'9R?�j�    IEND�B`�  THistoryComboBoxRemoteDirectoryEditLeft1TopTWidth�HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeControlChange  THistoryComboBoxLocalDirectoryEditLeft1Top#WidthBHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder TextLocalDirectoryEditOnChangeControlChange  TButtonLocalDirectoryBrowseButtonLeftzTop!WidthKHeightAnchorsakTopakRight Caption   Bl&äddra...TabOrderOnClickLocalDirectoryBrowseButtonClick   TButtonOkButtonLeft� Top�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft;Top�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder	  	TGroupBoxOptionsGroupLeftTop� Width/HeightICaption   Alternativ för synkroniseringTabOrder
DesignSize/I  	TCheckBoxSynchronizeDeleteCheckLeftTopWidth� HeightCaption&Ta bort filerTabOrder OnClickControlChange  	TCheckBoxSynchronizeSelectedOnlyCheckLeft� Top,Width� HeightAnchorsakLeftakTopakRight CaptionBara &valda filerTabOrderOnClickControlChange  	TCheckBoxSynchronizeExistingOnlyCheckLeft� TopWidth� HeightAnchorsakLeftakTopakRight Caption&Endast existerande filerTabOrderOnClickControlChange  	TCheckBoxSynchronizePreviewChangesCheckLeftTop,Width� HeightCaption   Fö&rhandsvisa ändringarTabOrderOnClickControlChange   TButtonTransferSettingsButtonLeftTop�Width� HeightAnchorsakLeftakBottom Caption   Överf&öringsinställningar...TabOrderOnClickTransferSettingsButtonClickOnDropDownClick#TransferSettingsButtonDropDownClick  	TGroupBoxDirectionGroupLeftTop� Width�Height1AnchorsakLeftakTopakRight Caption   Riktning/målkatalogTabOrder TRadioButtonSynchronizeBothButtonLeftTopWidth� HeightCaption   &BådaTabOrder OnClickControlChange  TRadioButtonSynchronizeRemoteButtonLeft� TopWidth� HeightCaption   &FjärrTabOrderOnClickControlChange  TRadioButtonSynchronizeLocalButtonLeft0TopWidth� HeightCaption&LokalTabOrderOnClickControlChange   	TGroupBoxCompareCriterionsGroupLeft=Top� Width� HeightIAnchorsakLeftakTopakRight Caption   JämförelsekriterierTabOrder
DesignSize� I  	TCheckBoxSynchronizeByTimeCheckLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption   Ä&ndringstidTabOrder OnClickControlChange  	TCheckBoxSynchronizeBySizeCheckLeftTop,Width� HeightAnchorsakLeftakTopakRight CaptionF&ilstorlekTabOrderOnClickControlChange   	TCheckBoxSaveSettingsCheckLeftTop=Width�HeightAnchorsakLeftakTopakRight Caption   Använd &samma val nästa gångTabOrder  	TGroupBoxCopyParamGroupLeftTopRWidth�Height2AnchorsakLeftakTopakRight Caption   ÖverföringsinställningarTabOrderOnClickCopyParamGroupClickOnContextPopupCopyParamGroupContextPopup
DesignSize�2  TLabelCopyParamLabelLeftTopWidth�HeightAnchorsakLeftakTopakRightakBottom AutoSizeCaptionCopyParamLabelWordWrap	OnClickCopyParamGroupClick   TButton
HelpButtonLeft�Top�WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrder
OnClickHelpButtonClick  	TGroupBox	ModeGroupLeftTop� Width�Height1AnchorsakLeftakTopakRight CaptionMetodTabOrder TRadioButtonSynchronizeFilesButtonLeftTopWidth� HeightCaptionSynkronisera &filerTabOrder OnClickControlChange  TRadioButtonMirrorFilesButtonLeft� TopWidth� HeightCaptionS&pegelfilerTabOrderOnClickControlChange  TRadioButtonSynchronizeTimestampsButtonLeft0TopWidth� HeightCaption   Synkronisera tidss&tämplarTabOrderOnClickControlChange    TPF0TImportSessionsDialogImportSessionsDialogLeftjTop� HelpType	htKeywordHelpKeyword	ui_importBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionImport sitesXClientHeightClientWidthwColor	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnShowFormShow
DesignSizew PixelsPerInch`
TextHeight TLabelLabelLeftTopWidth=HeightAnchorsakLeftakTopakRight Caption   &Importera från:  TButtonOKButtonLeft� Top� WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top� WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  	TListViewSessionListView2LeftTop#WidthiHeight� AnchorsakLeftakTopakRightakBottom 
Checkboxes	ColumnsWidth�   ColumnClickDoubleBuffered	HideSelectionReadOnly	ParentDoubleBufferedParentShowHintShowColumnHeadersShowHint	TabOrder	ViewStylevsReport	OnInfoTipSessionListView2InfoTipOnKeyUpSessionListView2KeyUpOnMouseDownSessionListView2MouseDown  TButtonCheckAllButtonLeftTop� WidthlHeightAnchorsakLeftakBottom CaptionMarkera/avmarkera &allaTabOrderOnClickCheckAllButtonClick  	TCheckBoxImportKeysCheckLeftTop� WidthYHeightAnchorsakLeftakBottom Caption4   Importera cachade &värdnycklar för valda sessionerTabOrder  TButton
HelpButtonLeft&Top� WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  	TComboBoxSourceComboBoxLeftjTopWidthxHeightStylecsDropDownListTabOrder OnSelectSourceComboBoxSelectItems.StringsPuTTY	Filezilla       TPF0TLicenseDialogLicenseDialogLeft�Top� ActiveControlCloseButtonBorderIconsbiSystemMenu BorderStylebsDialogCaption   AnvändarlicensClientHeight@ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenter
DesignSize�@ PixelsPerInch`
TextHeight TButtonCloseButtonLeft�TopWidthKHeightAnchorsakRightakBottom Cancel	Caption   StängDefault	ModalResultTabOrder   TMemoLicenseMemoLeftTopWidth�HeightAnchorsakLeftakTopakRight Color	clBtnFaceReadOnly	
ScrollBars
ssVerticalTabOrderWantReturns      TPF0TLocationProfilesDialogLocationProfilesDialogLeftWTop� HelpType	htKeywordHelpKeywordui_locationprofileBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionPlatsprofilerClientHeight�ClientWidth-Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnShowFormShow
DesignSize-� PixelsPerInch`
TextHeight TLabelLocalDirectoryLabelLeft.TopWidthJHeightCaptionL&okal katalog:FocusControlLocalDirectoryEdit  TLabelRemoteDirectoryLabelLeft.Top8WidthWHeightCaption   F&järrkatalog:FocusControlRemoteDirectoryEdit  TImageImageLeftTopWidth Height AutoSize	Picture.Data
*  	TPngImage�PNG

   IHDR           szz�   	pHYs  �  ��o�d  �IDATx��{L[Uǿ����e�.��X��P������l��F�4`��b��l#օ�(�m�_��h�7a5Ƃc�=�M�ɻ��aK�V�����ʥ��1����9���9����~���a4X#����#�=�j���]�3��J��M��� ���wLc��}�ɂ��ާJ��aY� �H�DkfS���Oh�' Q����8�P p��ÿ#nLx����
�^o��\7���ژ�'�Ts�t���
+Xe�����cN�ɉ۸��mR�������.��2>�}��(�O2h�����J�I�D�>��*NC��PA���vv׀�j�PO*+����&ĕV��g<רJ�Y�{������pc�Ht��8��z<k�Z��Sq�ĝە�t�Kj��J_<d,<,+?`�C������;/p<k�!����{��Q�Q��dDr:+;�h��,�)i�Ԋg_��q}�:^�Zz�i���eSX�j<�L��	~��˂�\�L���R7���������K-�w�F j�:�ʶfoڲa������%c� ����O��ܜ��+^\�Ͷ�( r�:o�5)ioX;q����}�l�͉G�eX4٬� �_2�
���hpN,�#"["x^�* ���S�sJ
_��ٹö�#ck�2��)L��� B��y�]��w��N�p�������$ ��C�x���ض�-`����G"��qԜϬ��yF&���y�:�/�Y `�&����`0e���)�T��X���1t�:NP�j	@IA� ��G����zH(�\�o��ˏ�NH ��׺���:��e�:u?�Pt?���3���+���H �41�ڣ��7���Nb���(�
-�(�8�mo(>�hJ-�i	@f�1���ʃ��5��"|,�CmD�tk�sC���f�� RX����,����y�;dQ��m��ƿ.�q���aa,ޅ�i*zܐ�ߜ��N�� ��}�CG�G�y���ďR�'�!�b�I�g�Z�=p��v��8~�`�ў�Jp�,��J�ZP#1����`��ː;
`���� N����Ő����� "~��"l�|N���y]	�f�	����Sr�hc�P*B"ZX�D$�sӅ?���w�Y k��d�=OB��b H�r�R���7(~@���T��:]jL�-��p}8�����Q���(��ڴa�k����a���V��j���FT��5�    IEND�B`�  TButtonOKBtnLeft/Top�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft�Top�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TPageControlPageControlLeftTophWidthHeight 
ActivePageSessionProfilesSheetAnchorsakLeftakTopakRightakBottom TabOrder 	TTabSheetSessionProfilesSheetTagCaptionSessionsplatsprofiler
DesignSize  	TTreeViewSessionProfilesViewTagLeft
Top	Width�Height� AnchorsakLeftakTopakRightakBottom DoubleBuffered	DragModedmAutomaticHideSelectionImagesBookmarkImageListIndentParentDoubleBufferedTabOrder OnChangeProfilesViewChangeOnCollapsedProfilesViewCollapsed
OnDblClickProfilesViewDblClick
OnDragDropProfilesViewDragDrop
OnDragOverProfilesViewDragOverOnEditedProfilesViewEdited	OnEditingProfilesViewEditing	OnEndDragProfilesViewEndDrag
OnExpandedProfilesViewExpandedOnGetImageIndexProfilesViewGetImageIndexOnGetSelectedIndexProfilesViewGetSelectedIndex	OnKeyDownProfilesViewKeyDownOnStartDragProfilesViewStartDragItems.NodeData
                ��������           1 "           ��������            1 1             ��������            2             ��������            3            ��������           4 "           ��������            4 1             ��������            5   TButtonAddSessionBookmarkButtonTagLeft�Top	WidthSHeightAnchorsakTopakRight Caption   &Lägg till...TabOrderOnClickAddBookmarkButtonClick  TButtonRemoveSessionBookmarkButtonTagLeft�Top)WidthSHeightAnchorsakTopakRight Caption&Ta bortTabOrderOnClickRemoveBookmarkButtonClick  TButtonDownSessionBookmarkButtonTagLeft�Top� WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickBookmarkButtonClick  TButtonUpSessionBookmarkButtonTag�Left�Top� WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickBookmarkButtonClick  TButtonRenameSessionBookmarkButtonTagLeft�TopIWidthSHeightAnchorsakTopakRight Caption	B&yt namnTabOrderOnClickRenameBookmarkButtonClick  TButtonSessionBookmarkMoveToButtonTagLeft�TopiWidthSHeightAnchorsakTopakRight Caption&Flytta till...TabOrderOnClickBookmarkMoveToButtonClick   	TTabSheetSharedProfilesSheetTagCaptionDelade platsprofiler
ImageIndex
DesignSize  	TTreeViewSharedProfilesViewTagLeft
Top	Width�Height� AnchorsakLeftakTopakRightakBottom DoubleBuffered	DragModedmAutomaticHideSelectionImagesBookmarkImageListIndentParentDoubleBufferedTabOrder OnChangeProfilesViewChangeOnCollapsedProfilesViewCollapsed
OnDblClickProfilesViewDblClick
OnDragDropProfilesViewDragDrop
OnDragOverProfilesViewDragOverOnEditedProfilesViewEdited	OnEditingProfilesViewEditing	OnEndDragProfilesViewEndDrag
OnExpandedProfilesViewExpandedOnGetImageIndexProfilesViewGetImageIndexOnGetSelectedIndexProfilesViewGetSelectedIndex	OnKeyDownProfilesViewKeyDownOnStartDragProfilesViewStartDragItems.NodeData
                ��������           1 "           ��������            1 1             ��������            2             ��������            3            ��������           4 "           ��������            4 1             ��������            5   TButtonAddSharedBookmarkButtonTagLeft�Top	WidthSHeightAnchorsakTopakRight Caption   &Lägg till...TabOrderOnClickAddBookmarkButtonClick  TButtonRemoveSharedBookmarkButtonTagLeft�Top)WidthSHeightAnchorsakTopakRight Caption&Ta bortTabOrderOnClickRemoveBookmarkButtonClick  TButtonRenameSharedBookmarkButtonTagLeft�TopIWidthSHeightAnchorsakTopakRight Caption	B&yt namnTabOrderOnClickRenameBookmarkButtonClick  TButtonSharedBookmarkMoveToButtonTagLeft�TopiWidthSHeightAnchorsakTopakRight Caption&Flytta till...TabOrderOnClickBookmarkMoveToButtonClick  TButtonUpSharedBookmarkButtonTag�Left�Top� WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickBookmarkButtonClick  TButtonDownSharedBookmarkButtonTagLeft�Top� WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickBookmarkButtonClick  TButtonShortCutSharedBookmarkButtonTagLeft�Top� WidthSHeightAnchorsakTopakRight Caption   &Genväg...TabOrderOnClickShortCutBookmarkButtonClick    TIEComboBoxLocalDirectoryEditLeft.TopWidth�HeightAnchorsakLeftakTopakRight TabOrder TextLocalDirectoryEditOnChangeDirectoryEditChange  TIEComboBoxRemoteDirectoryEditLeft.TopIWidth�HeightAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeDirectoryEditChange  TButtonLocalDirectoryBrowseButtonLeft�TopWidthKHeightAnchorsakTopakRight Caption   Blädd&ra...TabOrderOnClickLocalDirectoryBrowseButtonClick  TButtonSwitchButtonLeftTop�WidthaHeightAnchorsakRightakBottom Caption   &Bokmärken...ModalResultTabOrderOnClickSwitchButtonClick  TButton
HelpButtonLeft�Top�WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TPngImageListBookmarkImageList	PngImages
BackgroundclWindowNameBookmarkPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?%�����ɈEn?�m�&w�ܟG�@�3�xj�JK�b�P�����R?~�Ƹ�Y.DP�g���&��[�3�{�9����ƙ|����x$��~���p��i?	2nj��l�#$ƅb��W���f�|������.��l`����2 `���G��_W�_cp4���a�.����)�,��� lܾa�o��,V3c�SW�
�o�wɀ�T��ב��#(�[�a�U�f`g����)$2#~�Gр� ���l�Ԁ�@8uɀT/�?��l1�\`{��FJ���b��W�H�f`��I�+�.p8�`#"�����o�va���ÿ�X��?ܜ�Q�l%��	����a۝|R�Qm�b��)V���޽g0f���)܀O�4�7��2\����P�����O�ID  �/����>���I����ß?$�H)2��1|�r��~�d  m��7_��    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  iIDATx�c���?%�����ɈEn?�m�&w�ܟG�@�x��,"(ɿ�:� E���^|�y���Z�Z��h	I�H�{����+���yd3�k�6I�޽�*� F��	�$�y�y4�t.�|����;#��A��c�K�L�����3l�6@�L���Wms�?o����B#���G��0\:tw� Q	}5Q����©	�>����ǟ����13�j103~��-L!���20�X}�ǿ���HJr2���m�UȀd 
��~��p���~5=��9�0��)!�3��G�u���W3}k�`��,�(&BR�10|g��Oƣ��;F�s#�  6|�j���    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATx�c���?%�����ɈEn?�m�&w�ܟG�@��4�,f��,"(����GE��-�޽��W�x#^6��]��P��BQ���7��;�aw6�1���0���Ȓ���[3�V?d�@N��[y�$͛�M��Ne`�}9��J h���9'�Ȍ``�u�t�7�?�f@�ß���ۼ�2�����I�+��`�T����\�Q} ;t�%�>��N�j��e�>i^R��?��/~Տ�z)΍�  Tؚ�hƕ2    IEND�B`�  Left� Top�Bitmap
       TPF0TLogFormLogFormLeftdTop� HelpType	htKeywordHelpKeywordui_logBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp CaptionLogClientHeight/ClientWidth�Color	clBtnFaceConstraints.MinHeight� Constraints.MinWidth� 
ParentFont	OldCreateOrderOnClose	FormClosePixelsPerInch`
TextHeight TTBXStatusBar	StatusBarLeft TopWidth�HeightPanelsFramedMaxSize� Size� StretchPrioritydTag   UseSystemFont  TTBXDockTopDockLeft Top Width�Height	AllowDrag TTBXToolbarToolbarLeft Top CaptionToolbarFullSize	ImagesGlyphsModule.LogImagesParentShowHintShowHint	TabOrder  TTBXItemTBXItem2Action"NonVisualDataModule.LogClearAction  TTBXItemTBXItem3Action!NonVisualDataModule.LogCopyAction  TTBXItemTBXItem4Action&NonVisualDataModule.LogSelectAllAction  TTBXSeparatorItemTBXSeparatorItem2  TTBXItemTBXItem5Action(NonVisualDataModule.LogPreferencesAction        TPF0TLoginDialogLoginDialogLeft_Top� HelpType	htKeywordHelpKeywordui_loginBorderIconsbiSystemMenu
biMinimizebiHelp Caption
InloggningClientHeight�ClientWidthvColor	clBtnFaceConstraints.MinHeight^Constraints.MinWidthX
ParentFont	
KeyPreview	OldCreateOrder	PositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShowPixelsPerInch`
TextHeight TPanel	MainPanelLeftTop WidthiHeight�AlignalClient
BevelOuterbvNoneTabOrder  TPanelContentsPanelLeft Top WidthiHeight�AlignalClient
BevelOuterbvNoneTabOrder Visible
DesignSizei�  	TGroupBoxContentsGroupBoxLeftTopWidth[HeightxAnchorsakLeftakTopakBottom CaptionContentsGroupBoxTabOrder 
DesignSize[x  TLabelContentsLabelLeftTopWidthHeightCaptionNamn:  TEditContentsNameEditLeftBTopWidthHeightAnchorsakLeftakTopakRight TabOrder TextContentsNameEdit  TMemoContentsMemoLeftTop*WidthDHeightBAnchorsakLeftakTopakRightakBottom Lines.StringsContentsMemo TabOrder    TPanel	SitePanelLeft Top WidthiHeight�AlignalClientAnchorsakTopakRightakBottom 
BevelOuterbvNoneTabOrder
DesignSizei�  	TGroupBox
BasicGroupLeftTopWidth[Height� AnchorsakLeftakTopakRight CaptionSessionTabOrder 
DesignSize[�   TLabelLabel1LeftTopHWidth7HeightCaption   &Värdnamn:FocusControlHostNameEdit  TLabelLabel2Left� TopHWidth?HeightAnchorsakTopakRight CaptionPo&rtnummer:FocusControlPortNumberEdit  TLabelLabel3LeftTopzWidth7HeightCaption   &Användarnamn:FocusControlUserNameEdit  TLabelLabel4Left� TopzWidth2HeightCaption   &Lösenord:FocusControlPasswordEdit  TLabelLabel22LeftTopWidth>HeightCaption&Filprotokoll:FocusControlTransferProtocolCombo  TLabel	FtpsLabelLeft� TopWidth7HeightCaption&Kryptering:FocusControl	FtpsCombo  TLabelWebDavsLabelLeft� TopWidth7HeightCaption&Kryptering:FocusControlWebDavsCombo  TEditEncryptionViewLeft� Top'Width� HeightTabOrderOnChangeTransferProtocolComboChange  TEditTransferProtocolViewLeftTop'Width� HeightTabOrderOnChangeTransferProtocolComboChange  TEditHostNameEditLeftTopYWidth� HeightAnchorsakLeftakTopakRight 	MaxLengthdTabOrderTextHostNameEditOnChange
DataChange  TEditUserNameEditLeftTop� Width� Height	MaxLengthdTabOrderTextUserNameEditOnChange
DataChange  TPasswordEditPasswordEditLeft� Top� Width� HeightAnchorsakLeftakTopakRight 	MaxLengthdTabOrderTextPasswordEditOnChange
DataChange  TUpDownEditPortNumberEditLeft� TopYWidthRHeight	AlignmenttaRightJustifyMaxValue      ��@MinValue       ��?Value       ��?AnchorsakTopakRight TabOrderOnChangePortNumberEditChange  	TComboBoxTransferProtocolComboLeftTop'Width� HeightStylecsDropDownListTabOrder OnChangeTransferProtocolComboChangeItems.StringsSFTPSCPFTP   	TComboBox	FtpsComboLeft� Top'Width� HeightStylecsDropDownListTabOrderOnChangeTransferProtocolComboChangeItems.StringsIngen krypteringTLS/SSL Implicit encryptionXTLS Explicit encryptionXSSL Explicit encryptionX   	TComboBoxWebDavsComboLeft� Top'Width� HeightStylecsDropDownListTabOrderOnChangeTransferProtocolComboChangeItems.StringsNo encryptionXTLS/SSL Implicit encryptionX   TPanelBasicFtpPanelLeftTop� WidthDHeightAnchorsakLeftakTopakRight 
BevelOuterbvNoneTabOrder	 	TCheckBoxAnonymousLoginCheckLeft Top Width� HeightCaption&Anonym inloggningTabOrder OnClickAnonymousLoginCheckClick   TPanelBasicSshPanelLeftTop� Width[Height AnchorsakLeftakTopakRight 
BevelOuterbvNoneTabOrder
  TButtonAdvancedButtonLeft� Top� WidthbHeightActionSessionAdvancedActionAnchorsakRightakBottom StylebsSplitButtonTabOrderOnDropDownClickAdvancedButtonDropDownClick  TButton
SaveButtonLeftTop� Width`HeightActionSaveSessionActionAnchorsakLeftakBottom StylebsSplitButtonTabOrderOnDropDownClickSaveButtonDropDownClick  TButtonEditCancelButtonLefttTop� WidthRHeightActionEditCancelActionAnchorsakLeftakBottom TabOrderOnDropDownClickSaveButtonDropDownClick  TButton
EditButtonLeftTop� WidthbHeightActionEditSessionActionAnchorsakLeftakBottom TabOrderOnDropDownClickSaveButtonDropDownClick    TPanelButtonPanelLeft Top�WidthiHeight)AlignalBottom
BevelOuterbvNoneTabOrder
DesignSizei)  TButtonLoginButtonLeftKTop
WidthbHeightActionLoginActionAnchorsakRightakBottom Default	ImagesActionImageListModalResultStylebsSplitButtonTabOrder OnDropDownClickLoginButtonDropDownClick  TButtonCloseButtonLeft� Top
WidthRHeightAnchorsakRightakBottom Cancel	Caption   StängModalResultTabOrder  TButton
HelpButtonLeftTop
WidthRHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick    TPanel
SitesPanelLeft Top WidthHeight�AlignalLeftAnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneTabOrder
DesignSize�  	TTreeViewSessionTreeLeftTopWidth� HeightAnchorsakLeftakTopakRightakBottom DoubleBuffered	DragModedmAutomaticHideSelectionImagesSessionImageListIndentParentDoubleBufferedParentShowHint	RowSelect	ShowHint	ShowRootSortTypestBothTabOrder OnChangeSessionTreeChange
OnChangingSessionTreeChangingOnCollapsedSessionTreeExpandedCollapsed	OnCompareSessionTreeCompareOnContextPopupSessionTreeContextPopupOnCustomDrawItemSessionTreeCustomDrawItem
OnDblClickSessionTreeDblClick
OnDragDropSessionTreeDragDropOnEditedSessionTreeEdited	OnEditingSessionTreeEditing	OnEndDragSessionTreeEndDragOnExitSessionTreeExitOnExpandingSessionTreeExpanding
OnExpandedSessionTreeExpandedCollapsed	OnKeyDownSessionTreeKeyDown
OnKeyPressSessionTreeKeyPressOnMouseDownSessionTreeMouseDownOnMouseMoveSessionTreeMouseMoveOnStartDragSessionTreeStartDrag  TStaticTextSitesIncrementalSearchLabelLeftTopwWidth� HeightAnchorsakLeftakRightakBottom BorderStyle	sbsSingleCaptionSitesIncrementalSearchLabelShowAccelCharTabOrderVisible  TButtonManageButtonLeft� Top�WidthbHeightAnchorsakRightakBottom Caption&HanteraTabOrderOnClickManageButtonClick  TButtonToolsMenuButtonLeftTop�WidthbHeightAnchorsakLeftakBottom Caption&VerktygTabOrderOnClickToolsMenuButtonClick   TActionList
ActionListImagesActionImageListOnUpdateActionListUpdateLeftDTopQ TActionEditSessionActionCategorySessionsCaption	&Redigera	OnExecuteEditSessionActionExecute  TActionSaveAsSessionActionCategorySessionsCaption
&Spara somShortCutA�  	OnExecuteSaveAsSessionActionExecute  TActionSaveSessionActionCategorySessionsCaption	&Spara...	OnExecuteSaveSessionActionExecute  TActionDeleteSessionActionCategorySessionsCaptionTa &bort...
ImageIndex	OnExecuteDeleteSessionActionExecute  TActionImportSessionsActionCategorySessionsCaption&Importera...	OnExecuteImportSessionsActionExecute  TActionLoginActionCategorySessionCaptionLogga in
ImageIndex 	OnExecuteLoginActionExecute  TActionAboutActionCategoryOtherCaption&Om...	OnExecuteAboutActionExecute  TActionCleanUpActionCategoryOtherCaption&Rensa applikationsdata...	OnExecuteCleanUpActionExecute  TActionResetNewSessionActionCategorySessionsCaption   Å&terställ	OnExecuteResetNewSessionActionExecute  TActionSetDefaultSessionActionCategorySessionsCaption   Sä&tt som standard	OnExecuteSetDefaultSessionActionExecute  TActionDesktopIconActionCategorySessionsCaptionSkrivbords&ikon	OnExecuteDesktopIconActionExecute  TActionSendToHookActionCategorySessionsCaption"   Utforskarens 'Skicka till'-genväg	OnExecuteSendToHookActionExecute  TActionCheckForUpdatesActionTagCategoryOtherCaption   Sök efter &uppdateringar
ImageIndex?	OnExecuteCheckForUpdatesActionExecute  TActionRenameSessionActionCategorySessionsCaption	Byt &namn
ImageIndex	OnExecuteRenameSessionActionExecute  TActionNewSessionFolderActionCategorySessionsCaptionN&y katalog...
ImageIndex	OnExecuteNewSessionFolderActionExecute  TActionRunPageantActionCategoryOtherCaption   Kör &Pageant	OnExecuteRunPageantActionExecute  TActionRunPuttygenActionCategoryOtherCaption   Kör PuTTY&gen	OnExecuteRunPuttygenActionExecute  TActionImportActionCategoryOtherCaption'   Importera/Återställ &konfiguration...	OnExecuteImportActionExecute  TActionExportActionCategoryOtherCaption-   &Exportera/Säkerhetskopiera konfiguration...	OnExecuteExportActionExecute  TActionPreferencesActionCategoryOtherCaption   &Inställningar...	OnExecutePreferencesActionExecute  TActionEditCancelActionCategorySessionCaption&Avbryt	OnExecuteEditCancelActionExecute  TActionSessionAdvancedActionCategorySessionCaption&Avancerad...	OnExecuteSessionAdvancedActionExecute  TActionPreferencesLoggingActionCategoryOtherCaption&Loggning...	OnExecutePreferencesLoggingActionExecute  TActionCloneToNewSiteActionCategorySessionCaption&Klona till ny webbplats	OnExecuteCloneToNewSiteActionExecute  TActionPuttyActionCategorySessionCaption   Öppna i &PuTTY
ImageIndexShortCutP@SecondaryShortCuts.StringsShift+Ctrl+P 	OnExecutePuttyActionExecute   
TPopupMenuToolsPopupMenuLeft� Top�  	TMenuItemImport1ActionImportSessionsAction  	TMenuItemN3Caption-  	TMenuItemImportConfiguration1ActionImportAction  	TMenuItemExportConfiguration1ActionExportAction  	TMenuItemCleanup1ActionCleanUpAction  	TMenuItemN2Caption-  	TMenuItemPageant1ActionRunPageantAction  	TMenuItem	Puttygen1ActionRunPuttygenAction  	TMenuItemN1Caption-  	TMenuItemCheckForUpdates1ActionCheckForUpdatesAction  	TMenuItemN4Caption-  	TMenuItemPreferences1ActionPreferencesAction  	TMenuItemAbout1ActionAboutAction   TPngImageListSessionImageList	PngImages
BackgroundclWhiteNameUnusedPngImage.Data
b   �PNG

   IHDR         ��h6   tRNS �   ���/�   IDATx�c����8�aT���  �E�/UY"    IEND�B`� 
BackgroundclWindowNameSitePngImage.Data
J  �PNG

   IHDR         ��h6   tRNS � � �7X}   �IDATx�c���?)��d�IϞ�$�NJR|�� ��ދ������������P�?�rA��S�@5L��谿���p�.T��IC�� Q�:	R��d�1�:���5HHP��_�����������ן�����j���k�Ƽ��������T`z��(����������_(]���`���`����`�����C}d5jx|�TC`dʓg�I�i��d��gC�DOKp�J��6�S+ ����>�7    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  iIDATx�c���?%�����ɈEn?�m�&w�ܟG�@�x��,"(ɿ�:� E���^|�y���Z�Z��h	I�H�{����+���yd3�k�6I�޽�*� F��	�$�y�y4�t.�|����;#��A��c�K�L�����3l�6@�L���Wms�?o����B#���G��0\:tw� Q	}5Q����©	�>����ǟ����13�j103~��-L!���20�X}�ǿ���HJr2���m�UȀd 
��~��p���~5=��9�0��)!�3��G�u���W3}k�`��,�(&BR�10|g��Oƣ��;F�s#�  6|�j���    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATx�c���?%�����ɈEn?�m�&w�ܟG�@��4�,f��,"(����GE��-�޽��W�x#^6��]��P��BQ���7��;�aw6�1���0���Ȓ���[3�V?d�@N��[y�$͛�M��Ne`�}9��J h���9'�Ȍ``�u�t�7�?�f@�ß���ۼ�2�����I�+��`�T����\�Q} ;t�%�>��N�j��e�>i^R��?��/~Տ�z)΍�  Tؚ�hƕ2    IEND�B`� 
BackgroundclWindowName	WorkspacePngImage.Data
/  �PNG

   IHDR         ��h6   tRNS � � �7X}   �IDATx�c���?)��d�A-���!F���ȥ�Ռ<f���h8�����~�������Ԁ�0oѪ��0	��Ahx~�Ͱ����m�%�J����t�P��J� �-K���ؠ	�9�B5��ӅfX����h�J.eP7wv�8u(�a�d ��UǊì���ˡ�l�@3l���y��h�:^P�7���M�p"3�M�з�!-ٟ�x�5w#NOcPO���HM� WՌ�\[    IEND�B`� 
BackgroundclWindowNameWorkspace closedPngImage.Data
b   �PNG

   IHDR         ��h6   tRNS �   ���/�   IDATx�c����8�aT���  �E�/UY"    IEND�B`� 
BackgroundclWindowNameNew Site openedPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�cd ���``d���)��!�WL�Lɟ?���͸�H����d��>����7Y��~��[��+����89�l��׷��fx����/�=xe��+�^��g�����3T�c���c�d����쵇N_�߸�+������P�"6ظ���M|����M8�X��g`�}������z�d��)��%�3 ���H��d��w>3�>w�!�ǂAJT��ś��w�e�q������OY���1�ç��Na�a`fbb��g�u��敝�~ W���_�5 �f`x��1ã�w�5~���p���?��Vv��(�^������>1����?÷_@��l�b�ѵ�^љvn@^����|���������3���=f.�f8}p+<���6lfx����M���$_L��� ���DLd5�6������D���ph�� l*@����m�qiD� :�lV�B    IEND�B`� 
BackgroundclWindowNameNew Site closedPngImage.Data
r   �PNG

   IHDR         ��h6   sRGB ���   	pHYs  �  ��o�d   IDATx�c���?)�qTè�� ��/�Ǭ�Y    IEND�B`� 
BackgroundclWindowNameSite color maskPngImage.Data
�   �PNG

   IHDR         ��h6   tRNS � � �@�   bIDATx�c�����H����g�_T'%)��pH���w��K54D��:<���d5jx|�TC`dʓg�	j@�4ZZ2+���!F��d�� Mɩ �ROqe�!�    IEND�B`�  LeftDTopBitmap
      
TPopupMenuSaveDropDownMenuLeftDTop�  	TMenuItemSaveSessionMenuItemActionSaveSessionActionDefault	  	TMenuItemSaveAsSessionMenuItemActionSaveAsSessionAction  	TMenuItemN7Caption-  	TMenuItemSetdefaults1ActionSetDefaultSessionAction   
TPopupMenuManageSitePopupMenuImagesActionImageListLeftDTop�  	TMenuItem
Shellicon1Caption	WebbplatsEnabledVisible  	TMenuItemSiteLoginMenuItemActionLoginActionDefault	  	TMenuItemOpeninPuTTY2ActionPuttyAction  	TMenuItemN10Caption-  	TMenuItemEdit1ActionEditSessionAction  	TMenuItemDelete1ActionDeleteSessionAction  	TMenuItemRename1ActionRenameSessionAction  	TMenuItemSiteClonetoNewSiteMenuItemActionCloneToNewSiteAction  	TMenuItemN5Caption-  	TMenuItemSetdefaults2ActionSetDefaultSessionAction  	TMenuItemN6Caption-  	TMenuItem
Newfolder1ActionNewSessionFolderAction  	TMenuItem
Shellicon2CaptionIkon webbplatsEnabledVisible  	TMenuItemDesktopIcon2ActionDesktopIconAction  	TMenuItemExplorersSendToShortcut2ActionSendToHookAction   
TPopupMenuManageFolderPopupMenuImagesActionImageListLeftFTop	 	TMenuItem	MenuItem1CaptionWebbplatskatalogEnabledVisible  	TMenuItemLogin5ActionLoginActionDefault	  	TMenuItemN11Caption-  	TMenuItem	MenuItem3ActionDeleteSessionAction  	TMenuItem	MenuItem4ActionRenameSessionAction  	TMenuItem	MenuItem5Caption-  	TMenuItem	MenuItem6ActionNewSessionFolderAction  	TMenuItem	MenuItem7CaptionIkon webbplatskatalogEnabledVisible  	TMenuItem	MenuItem8ActionDesktopIconAction   
TPopupMenuManageNewSitePopupMenuImagesActionImageListLeft� Top�  	TMenuItem
MenuItem12CaptionNy webbplatsEnabledVisible  	TMenuItemLogin2ActionLoginActionDefault	  	TMenuItemOpeninPuTTY3ActionPuttyAction  	TMenuItemN8Caption-  	TMenuItem
MenuItem13ActionSaveAsSessionAction  	TMenuItemReset1ActionResetNewSessionAction  	TMenuItem
MenuItem21Caption-  	TMenuItem
MenuItem22ActionSetDefaultSessionAction  	TMenuItem
MenuItem16Caption-  	TMenuItem
MenuItem17ActionNewSessionFolderAction   
TPopupMenuManageWorkspacePopupMenuImagesActionImageListLeft� Top 	TMenuItem	MenuItem2Caption	ArbetsytaEnabledVisible  	TMenuItemLogin3ActionLoginActionDefault	  	TMenuItemN9Caption-  	TMenuItem
MenuItem10ActionDeleteSessionAction  	TMenuItem
MenuItem11ActionRenameSessionAction  	TMenuItem
MenuItem18CaptionIkon arbetsytaEnabledVisible  	TMenuItem
MenuItem19ActionDesktopIconAction   
TPopupMenuSessionAdvancedPopupMenuLeft� TopY 	TMenuItemSession1CaptionSessionEnabledVisible  	TMenuItem	MenuItem9ActionSessionAdvancedActionDefault	  	TMenuItem
MenuItem14Caption   Globala inställningarEnabledVisible  	TMenuItemPreferencesLoggingAction1ActionPreferencesLoggingAction   TPngImageListActionImageList	PngImages
BackgroundclWindowNameLoginPngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��o�d  �IDATx�cTh��!������ ���g*�|��oIavfR�3���������.�/�/\㰗A�S���ߟ0�p��]|� 6 ���1�[V[������⚂`��w,6����F=]������b �����CU �
��`�N�~��C����/�@V�������N=zL����a��.���3���,n�Z	,���G����"�����jO2�	<�`�\,���g�2<�c��gj�2�9�`�D,����|��.�?�{a�����炽 �_(����+� 1N���'��d��ǟ2��f����`d5_^}��%�����A{�4���8���H÷�_Q\���ۻ8����3�3hN���j~|�1���,�'���^�|z�������783��3�0222��������_pf�(; 1bҩCo��    IEND�B`� 
BackgroundclWindowNameOpen current session in PuTTYPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATxڅ�]HSa�g�meVt��6J�����.�0��""
��� �nv�]bA݈�1�>�"��8��bj�)i���)��R��<����ak{�����=���#��Qy`H��GP����XPAQ��G�M��.�%+�r��x�:"�Ǎ&/���;�����Of��7b���%n,%*���Dbs�����'(��c�f�>��,|��zMg��̀��2ŵ���1�������AL^�׵�D��lK�fY��3;��ؿ�$3�~���)Z'v�
?�)n���c�F��܀$�]���f&g��� O�-���������^!e��sa4ф���O��I�n����p[E�|���,TK�*/�*K�Ect>����(��k�W�F�cI��~�شX?
uW�����P�Z�f?O{c.������f](���̿��n���K��+<���'f���ׅ#�J�|�5����ʸ�� �"�Mg�)��01%�X���L6)WH������5�(�    IEND�B`� 
BackgroundclWindowNameRenamePngImage.Data
y  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�cd ���+-+���ɋ�'>,`$Es������'�uT����p��`�Ḫ\���`����:?���G�h6����h������_��'6nk��v~+��^�w��Z����GW�}[� F�@C����"g��op�����������y�$G�痛�Է2P���5ÍK7�m�U����Qln�p
�Z�)`��������W?�
�g/���fF���&��l���y�p��%�E�QՀXؒ�ՀgW�2Hrng`�Nexz���U��A@�._3b���$���yF���?d �A��5-1v��^�aP�bH؀���`����06\Z�ɠ������YQ�(nQ@��L�I �,`��A`Ru:���&��e(��4�A���U�3�/d�U�c�|��5�1e-�|��X��l@gY1��w-���  �����i�    IEND�B`� 
BackgroundclWindowNameDelete filePngImage.Data
z  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڥ�]HSaǟ�M�9�۔�t�ϴYJhe H!E7xQN*���Oꦫ��i	]TDA�`XMLYY:�3C��<�̹������$Q���}���<����B�'�� p��S!�nPO���V���|�J����=*I^��qN��^g�F˸ϯ,�m���wq'�Y���vǆ��	<C�vAr� �����RU�(.��b��y�D"��C����ss�4E�*/�;����y���/���7��YL��7WI HQx�i8�Jɻ	���Tߦ�{����&atb꣬��:67U	���\���﨩��`^����H��k+J,vk>��g�;��f�$�T��"^ m<{���9�XUM������d��0�O�irE"���V �����Z���3�lO��O�H ���X6w ��Ȼ��6ڨשg��2��7eF_���'t4yc���dqw!���͌Z�G�,^��`0�
p�gϲ4}��X�E\�e���4Bɭ�3�x�&S�X�Q��H.�F�*GQgx��8�AT�
j�m|����c��+��L>������5�|�^o2�TbK���S.Q���m$���i-6���Lɝح �V
��:�fF�i�\���VX�`(�~]I�v�4 �a�D�X�V,�}�{�%J���L]&}������T��Zp�7����x �D����LB����k�RFfP    IEND�B`� 
BackgroundclWindowNameCreate directoryPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�cd ���bd`���z�����/�j���?,|���o2c@X٬Yq����|<�����,,L�~��Zѝ������d�"���Mߑs�_�0�����n}>n�w�1�x������+�2�0nn���Ym�������&�d�72Ԑg���e�d���;ì��N_{X��+��qS��Uk%-!1.޽�ưi���B,̬��M�YY��g`�q�
�������d�WY���A�a��$�XosIQ��?0��}������1�_6 _ ~�+�p���AD������AB������=m�� �[y�G/<a8t����
��o?l� �wCu�R$�S~_G�����Rw^�2�x�!��8����cՀC�y�Y��GH�z10�y���?��P�͋.��h����#�dW`q����9+00���%��� *v��KT|R�1���c˜9(|Ҽ$������<�a���?)z1  �O�ہZ�    IEND�B`�  Left� TopBitmap
      
TPopupMenuLoginDropDownMenuImagesActionImageListLeftFTopA 	TMenuItemLogin1ActionLoginActionDefault	  	TMenuItemOpeninPuTTY1ActionPuttyAction      TPF0TNonVisualDataModuleNonVisualDataModuleOldCreateOrderHeight�Widthp TActionList
LogActionsImagesGlyphsModule.LogImages	OnExecuteLogActionsExecuteOnUpdateLogActionsUpdateLeft Toph TActionLogClearActionCategoryLogMemoCaption&RensaHint
Rensa logg
ImageIndex ShortCut.@  TActionLogSelectAllActionCategoryLogMemoCaptionM&arkera alltHintMarkera allt
ImageIndexShortCutA@  TActionLogCopyActionCategoryLogMemoCaption&KopieraHintKopiera till urklipp
ImageIndexShortCutC@  TActionLogPreferencesActionCategoryLogFormCaptionLogPreferencesActionHintKonfigurera loggning
ImageIndex   TTBXPopupMenuLogMemoPopupImagesGlyphsModule.LogImagesLeft Top�  TTBXItemClear1ActionLogClearAction  TTBXItemClose1ActionLogCopyAction  TTBXItem
Selectall1ActionLogSelectAllAction   TTBXPopupMenuRemoteFilePopupImagesGlyphsModule.ExplorerImagesLeft�TopP TTBXItem	TBXItem23ActionCurrentAddEditLinkContextAction  TTBXItemRemoteOpenMenuItemActionCurrentOpenAction  TTBXItemRemoteEditMenuItemActionCurrentEditFocusedAction  TTBXItemRemoteCopyMenuItemActionRemoteCopyFocusedAction  TTBXItemMoveto1ActionRemoteMoveFocusedAction  TTBXItem
Duplicate3ActionRemoteCopyToAction  TTBXItemMoveto6ActionRemoteMoveToFocusedAction  TTBXItemDelete1ActionCurrentDeleteFocusedAction  TTBXItemRename1ActionCurrentRenameAction  TTBXSeparatorItemN45  TTBXSubmenuItemRemoteDirViewCustomCommandsMenuActionCustomCommandsAction TTBXItem    TTBXSubmenuItem
FileNames3Caption&FilnamnHelpKeyword	filenamesHint$   Operationer med namn på valda filer TTBXItemInserttoCommandLine2ActionFileListToCommandLineAction  TTBXItemCopytoClipboard3ActionFileListToClipboardAction  TTBXItemCopytoClipboardIncludePaths3ActionFullFileListToClipboardAction  TTBXItemCopyURLtoClipboard3ActionUrlToClipboardAction   TTBXSeparatorItemN1  TTBXItemProperties1ActionCurrentPropertiesFocusedAction   TActionListExplorerActionsImagesGlyphsModule.ExplorerImages	OnExecuteExplorerActionsExecuteOnUpdateExplorerActionsUpdateLeft�Top TActionLocalCopyFocusedActionTagCategoryLocal Focused OperationCaption   &Överför...HelpKeywordtask_uploadHint3   Överför|Överför lokala filer till fjärrkatalog
ImageIndexX  TActionRemoteCopyFocusedActionTagCategoryRemote Focused OperationCaption&Ladda ner...HelpKeywordtask_downloadHint9   Ladda ner|Ladda ner fjärrfiler till den lokala katalogen
ImageIndexY  TActionRemoteMoveFocusedActionTagCategoryRemote Focused OperationCaptionLadda ner och &ta bort...HelpKeywordtask_downloadHint\   Ladda ner och ta bort|Ladda ner fjärrfiler till den lokala katalogen och ta bort originalet
ImageIndexa  TActionRemoteCopyActionTagCategoryRemote Selected OperationCaptionLadda &ner...HelpKeywordtask_downloadHint9   Ladda ner|Ladda ner fjärrfiler till den lokala katalogen
ImageIndexY  TActionBestFitColumnActionTagCategoryColumnsCaption   &Bästa passningHint6   Bästa passning|Anpassa kolumnbredden till innehållet  TActionGoToTreeActionTagCategoryViewCaption   Gå till trädHelpKeywordui_file_panel#directory_treeHint   Gå till träd
ImageIndexLShortCutT�    TActionLocalTreeActionTagCategoryViewCaption   &TrädHelpKeywordui_file_panel#directory_treeHint   Dölj/visa katalogträd
ImageIndexLShortCutT�    TActionRemoteTreeActionTagCategoryViewCaption   &TrädHelpKeywordui_file_panel#directory_treeHint   Dölj/visa katalogträd
ImageIndexLShortCutT�    TActionQueueItemQueryActionTagCategoryQueueCaption   Vi&sa frågaHelpKeywordui_queue#managing_the_queueHint'   Visa avvaktande fråga på vald köpost
ImageIndexC  TActionQueueItemErrorActionTagCategoryQueueCaption	Vi&sa felHelpKeywordui_queue#managing_the_queueHint.   Visa avvaktande felmeddelande på vald köpost
ImageIndexD  TActionQueueItemPromptActionTagCategoryQueueCaptionVi&sa promptHelpKeywordui_queue#managing_the_queueHint'   Visa avvaktande prompt på vald köpost
ImageIndexE  TActionGoToCommandLineActionTagCategoryViewCaption   Gå till komma&ndoradHelpKeywordui_commander#command_lineHint   Gå till kommandoradShortCutN`  TActionQueueItemDeleteActionTagCategoryQueueCaption&AvbrytHelpKeywordui_queue#managing_the_queueHint   Ta bort vald köpost
ImageIndexG  TActionQueueItemExecuteActionTagCategoryQueueCaption
   &Utför nuHelpKeywordui_queue#managing_the_queueHintC   Utför vald köpost omedelbart genom att ge den en extra anslutning
ImageIndexF  TActionSelectOneActionTagCategory	SelectionCaption&Markera/avmarkeraHelpKeywordui_file_panel#selecting_filesHint"Markera|Markera/avmarkera vald fil  TActionCurrentRenameActionTagCategorySelected OperationCaption	&Byt namnHelpKeywordtask_renameHint   Byt namn|Byt namn på vald fil
ImageIndex  TActionLocalSortAscendingActionTag	CategorySortCaption	Stig&andeHelpKeywordui_file_panel#sorting_filesHintT   Stigande/fallande|Växla mellan stigande och fallande sortering i den lokala panelen
ImageIndex%  TActionCurrentEditActionTagCategorySelected OperationCaption	&RedigeraHelpKeyword	task_editHintRedigera|Redigera markerad fil
ImageIndex9  TActionHideColumnActionTagCategoryColumnsCaption   &Dölj kolumnHelpKeywordui_file_panel#selecting_columnsHint   Dölj kolumn|Dölj vald kolumn  TActionLocalBackActionTag	CategoryLocal DirectoryCaption	Till&bakaHelpKeywordtask_navigate#special_commands
ImageIndexShortCut%�    TActionCurrentCycleStyleActionTagCategoryStyleCaptionVisaHelpKeywordui_file_panel#view_styleHint9   Visa|Växla mellan att visa olika stilar för katalogvyer
ImageIndex  TActionCurrentIconActionTagCategoryStyleCaptionSt&ora ikonerHelpKeywordui_file_panel#view_styleHintStora ikoner|Visa stora ikoner
ImageIndex  TActionCurrentSmallIconActionTagCategoryStyleCaption   &Små ikonerHelpKeywordui_file_panel#view_styleHint   Små ikoner|Visa små ikoner
ImageIndex	  TActionCurrentListActionTagCategoryStyleCaptionLis&taHelpKeywordui_file_panel#view_styleHintLista|Visa lista
ImageIndex
  TActionCurrentReportActionTagCategoryStyleCaption&Detaljerad listaHelpKeywordui_file_panel#view_styleHint&Detaljerad lista|Visa detaljerad lista
ImageIndex  TActionRemoteMoveToActionTagCategoryRemote Selected OperationCaption&Flytta till...HelpKeyword'task_move_duplicate#moving_remote_filesHint0   Flytta|Flytta markerade filer till fjärrkatalog
ImageIndexd  TActionCurrentDeleteFocusedActionTagCategoryFocused OperationCaption&Ta bortHelpKeywordtask_deleteHintTa bort|Ta bort markerade filer
ImageIndex  TActionCurrentPropertiesFocusedActionTagCategoryFocused OperationCaption&EgenskaperHelpKeywordtask_propertiesHint6   Egenskaper|Visa/ändra egenskaper för markerade filer
ImageIndex  TActionCurrentCreateDirActionTagCategorySelected OperationCaptionS&kapa katalog...HelpKeywordtask_create_directoryHintSkapa katalog|Skapa ny katalog
ImageIndex  TActionCurrentDeleteActionTagCategorySelected OperationCaption&Ta bortHelpKeywordtask_deleteHintTa bort|Ta bort markerade filer
ImageIndex  TActionCurrentPropertiesActionTagCategorySelected OperationCaption&EgenskaperHelpKeywordtask_propertiesHint6   Egenskaper|Visa/ändra egenskaper för markerade filer
ImageIndex  TActionRemoteBackActionTagCategoryRemote DirectoryCaption	Till&bakaHelpKeywordtask_navigate#special_commands
ImageIndexShortCut%�    TActionRemoteForwardActionTagCategoryRemote DirectoryCaption   &FramåtHelpKeywordtask_navigate#special_commands
ImageIndexShortCut'�    TActionCommandLinePanelActionTagCategoryViewCaptionKomma&ndoradHelpKeywordui_commander#command_lineHint   Dölj/visa kommandoradShortCutN`  TActionRemoteParentDirActionTagCategoryRemote DirectoryCaption   &Överliggande katalogHelpKeywordtask_navigate#special_commandsHint"   Huvudkatalog|Gå till huvudkatalog
ImageIndex  TActionRemoteRootDirActionTagCategoryRemote DirectoryCaption&RotkatalogHelpKeywordtask_navigate#special_commandsHint   Rotkatalog|Gå till rotkatalog
ImageIndexShortCut�@  TActionRemoteHomeDirActionTagCategoryRemote DirectoryCaption&HemkatalogHelpKeywordtask_navigate#special_commandsHint   Hemkatalog|Gå till hemkatalog
ImageIndex  TActionRemoteRefreshActionTagCategoryRemote DirectoryCaption
&UppdateraHint$   Uppdatera|Uppdatera kataloginnehåll
ImageIndex  TActionAboutActionTagCategoryHelpCaption&Om...HelpKeywordui_aboutHintOm|Visa programinformation
ImageIndexA  TActionStatusBarActionTagCategoryViewCaption   &StatusfältHint   Visa/dölj statusfältet  TActionSessionsTabsActionTagCategoryViewCaptionSessionsflikarHint   Dölj/visa sessionsflikar  TActionExplorerAddressBandActionTagCategoryViewCaption&AdressHelpKeywordui_toolbarsHint   Visa/dölj adressfältet  TActionExplorerMenuBandActionTagCategoryViewCaption&MenyHelpKeywordui_toolbarsHint   Visa/dölj meny  TActionExplorerToolbarBandActionTagCategoryViewCaption&StandardknapparHelpKeywordui_toolbarsHint"   Visa/dölj standardverktygsfältet  TActionRemoteOpenDirActionTagCategoryRemote DirectoryCaption   &Öppna katalog/bokmärkeHelpKeyword$task_navigate#entering_path_manuallyHintC   Öppna katalog/bokmärke|Öppna vald katalog eller sparat bokmärke
ImageIndex  TActionSelectActionTagCategory	SelectionCaption&Markera filerHelpKeyword	ui_selectHint Markera|Markera filer efter mask
ImageIndex  TActionUnselectActionTagCategory	SelectionCaptionA&vmarkera filerHelpKeyword	ui_selectHint$Avmarkera|Avmarkera filer efter mask
ImageIndex  TActionSelectAllActionTagCategory	SelectionCaptionM&arkera allaHelpKeywordui_file_panel#selecting_filesHintMarkera alla
ImageIndex  TActionInvertSelectionActionTagCategory	SelectionCaption&Invertera markeringHelpKeywordui_file_panel#selecting_filesHintInvertera markering
ImageIndex  TActionExplorerSelectionBandActionTagCategoryViewCaption&MarkeringsknapparHelpKeywordui_toolbarsHint)   Dölj/visa verktygsfältet för markering  TActionClearSelectionActionTagCategory	SelectionCaption&Rensa markeringHelpKeywordui_file_panel#selecting_filesHintRensa markering
ImageIndex  TActionExplorerSessionBandActionTagCategoryViewCaptionSessio&nsknapparHelpKeywordui_toolbarsHint)   Dölj/visa verktygsfältet för sessioner  TActionExplorerPreferencesBandActionTagCategoryViewCaption   InställningsknapparHelpKeywordui_toolbarsHint.   Visa/dölj verktygsfältet för inställningar  TActionExplorerSortBandActionTagCategoryViewCaptionSo&rteringsknapparHelpKeywordui_toolbarsHint)   Visa/dölj verktygsfältet för sortering  TActionExplorerUpdatesBandActionTagCategoryViewCaption&UppdateringsknappHelpKeywordui_toolbarsHint+   Dölj/visa verktygsfält för uppdateringar  TActionExplorerTransferBandActionTagCategoryViewCaption   &Överför inställningarHelpKeywordui_toolbarsHint9   Dölj/visa verktygsfält för överföringsinställningar  TAction ExplorerCustomCommandsBandActionTagCategoryViewCaptionEgna ko&mmandoknapparHelpKeywordui_toolbarsHint,   Dölj/visa verktygsfält för egna kommandon  TActionViewLogActionTagCategoryViewCaption   Lo&ggfönsterHelpKeywordui_logHint   Visa/dölj loggfönster
ImageIndex  TActionNewSessionActionTagCategorySessionCaption&Ny session...HelpKeyword.task_connections#opening_additional_connectionHintW   Ny session|Öppna ny session (Håll nere SHIFT för att öppna den i ett nytt fönster)
ImageIndexShortCutN@SecondaryShortCuts.StringsCtrl+Shift+N   TActionSiteManagerActionTagCategorySessionCaption&Hantera webbplats...HelpKeywordui_login_stored_sessionsHints   Hantera webbplats|Öppnar hantera webbplats (håll ner Shift för att öppna hantera webbplats i ett nytt fönster)  TActionCloseSessionActionTagCategorySessionCaption   &Koppla ifrånHint&   Stäng session|Avsluta aktuell session
ImageIndexShortCutD`SecondaryShortCuts.StringsCtrl+W   TActionSavedSessionsAction2TagCategorySessionCaptionWebb&platserHelpKeyword.task_connections#opening_additional_connectionHint   Öppna webbplats
ImageIndex  TActionWorkspacesActionTagCategorySessionCaption&ArbetsytorHelpKeyword	workspaceHint   Öppna arbetsyta
ImageIndexe  TActionPreferencesActionTagCategoryViewCaption   &Inställningar...HelpKeywordui_preferencesHint2   Inställningar|Visa/ändra användarinställningar
ImageIndexShortCutP�    TActionRemoteChangePathActionTagCategoryRemote DirectoryCaption&Byt katalogHelpKeywordtask_navigateHint1   Tillåter att annan katalog välj i fjärrpanelen
ImageIndexShortCutq�    TActionLocalForwardActionTag	CategoryLocal DirectoryCaption   &FramåtHelpKeywordtask_navigate#special_commands
ImageIndexShortCut'�    TActionLocalParentDirActionTagCategoryLocal DirectoryCaption&HuvudkatalogHelpKeywordtask_navigate#special_commandsHint"   Huvudkatalog|Gå till huvudkatalog
ImageIndex  TActionLocalRootDirActionTagCategoryLocal DirectoryCaption&RotkatalogHelpKeywordtask_navigate#special_commandsHint    Rotkatalog|Gå till rotkatalogen
ImageIndexShortCut�@  TActionLocalHomeDirActionTag	CategoryLocal DirectoryCaption&HemkatalogHelpKeywordtask_navigate#special_commandsHint    Hemkatalog|Gå till hemkatalogen
ImageIndex  TActionLocalRefreshActionTag	CategoryLocal DirectoryCaption
&UppdateraHint$   Uppdatera|Uppdatera kataloginnehåll
ImageIndex  TActionLocalOpenDirActionTag	CategoryLocal DirectoryCaption   &Öppna katalog/bokmärke...HelpKeyword$task_navigate#entering_path_manuallyHintC   Öppna katalog/bokmärke|Öppna vald katalog eller sparat bokmärke
ImageIndex  TActionLocalChangePathActionTagCategoryLocal DirectoryCaption
&Byt enhetHelpKeywordtask_navigateHint1   Tillåter att annan enhet väljs för lokal panel
ImageIndexShortCutp�    TActionToolBar2ActionTagCategoryViewCaption   Verktygsfält snabb&tangenterHelpKeywordui_toolbarsHint.   Dölj/visa verktygsfältet för snabbtangenter  TActionCommanderMenuBandActionTagCategoryViewCaption&MenyHelpKeywordui_toolbarsHint   Dölj/visa meny  TActionCommanderSessionBandActionTagCategoryViewCaptionSessio&nsknapparHelpKeywordui_toolbarsHint)   Dölj/visa verktygsfältet för sessioner  TActionCommanderPreferencesBandActionTagCategoryViewCaption   InställningsknapparHelpKeywordui_toolbarsHint.   Dölj/visa verktygsfältet för inställningar  TActionCommanderSortBandActionTagCategoryViewCaptionS&orteringsknapparHelpKeywordui_toolbarsHint)   Dölj/visa verktygsfältet för sortering  TActionCommanderUpdatesBandActionTagCategoryViewCaption&UppdateringsknappHelpKeywordui_toolbarsHint)   Dölj/visa verktygsfält för uppdatering  TActionCommanderTransferBandActionTagCategoryViewCaption   ÖverföringsinställningarHelpKeywordui_toolbarsHint9   Dölj/visa verktygsfält för överföringsinställningar  TActionCommanderCommandsBandActionTagCategoryViewCaption&KommandoknapparHelpKeywordui_toolbarsHint)   Visa/dölj verktygsfältet för kommandon  TAction!CommanderCustomCommandsBandActionTagCategoryViewCaptionEgna ko&mmandoknapparHelpKeywordui_toolbarsHint,   Dölj/visa verktygsfält för egna kommandon  TActionCommanderLocalHistoryBandActionTagCategoryViewCaption&HistorikknapparHelpKeywordui_toolbarsHint.   Dölj/visa verktygsfältet för lokal historik  TAction"CommanderLocalNavigationBandActionTagCategoryViewCaption&NavigeringsknapparHelpKeywordui_toolbarsHint0   Dölj/visa verktygsfältet för lokal navigering  TActionCommanderLocalFileBandActionTagCategoryViewCaption&FilknapparHelpKeywordui_toolbarsHint,   Dölj/visa verktygsfältet för lokala filer  TAction!CommanderLocalSelectionBandActionTagCategoryViewCaption&MarkeringsknapparHelpKeywordui_toolbarsHint6   Dölj/visa verktygsfält för lokala markeringsknappar  TAction CommanderRemoteHistoryBandActionTagCategoryViewCaption&HistorikknapparHelpKeywordui_toolbarsHint)   Dölj/visa verktygsfältet fjärrhistorik  TAction#CommanderRemoteNavigationBandActionTagCategoryViewCaption&NavigeringsknapparHelpKeywordui_toolbarsHint0   Dölj/visa verktygsfältet för fjärrnavigering  TActionCommanderRemoteFileBandActionTagCategoryViewCaption&FilknapparHelpKeywordui_toolbarsHint+   Dölj/visa verktygsfältet för fjärrfiler  TAction"CommanderRemoteSelectionBandActionTagCategoryViewCaption&MarkeringsknapparHelpKeywordui_toolbarsHint7   Visa/dölj verktygsfältet för fjärrmarkeringsknappar  TActionLocalStatusBarActionTagCategoryViewCaption   Statusf&ältHint*   Dölj/visa den lokala panelens statusfält  TActionRemoteStatusBarActionTagCategoryViewCaption   Statusf&ältHint%   Dölj/visa fjärrpanelens statusfält  TActionLocalSortByNameActionTag	CategorySortCaptionEfter &namnHelpKeywordui_file_panel#sorting_filesHint8Sortera efter namn|Sortera den lokala panelen efter namn
ImageIndexShortCutr@  TActionLocalSortByExtActionTag	CategorySortCaption   Efter &filändelseHelpKeywordui_file_panel#sorting_filesHintF   Sortera efter filändelse|Sortera den lokala panelen efter filändelse
ImageIndex ShortCuts@  TActionLocalSortBySizeActionTag	CategorySortCaptionEfter &storlekHelpKeywordui_file_panel#sorting_filesHintASortera efter storlek|Sortera den lokala panelen efter filstorlek
ImageIndex#ShortCutu@  TActionLocalSortByAttrActionTag	CategorySortCaptionEfter &attributHelpKeywordui_file_panel#sorting_filesHint@Sortera efter attribut|Sortera den lokala panelen efter attribut
ImageIndex$ShortCutv@  TActionLocalSortByTypeActionTag	CategorySortCaptionEfter fil&typHelpKeywordui_file_panel#sorting_filesHint<Sortera efter filtyp|Sortera den lokala panelen efter filtyp
ImageIndex"  TActionLocalSortByChangedActionTag	CategorySortCaption   Efter senast &ändradHelpKeywordui_file_panel#sorting_filesHintM   Sortera efter senast &ändrad|Sortera den lokala panelen efter senast ändrad
ImageIndex!ShortCutt@  TActionRemoteSortAscendingActionTagCategorySortCaption	Stig&andeHelpKeywordui_file_panel#sorting_filesHintW   Stigande/fallande|Växla sortering mellan stigande och fallande ordning i fjärrpanelen
ImageIndex%  TActionRemoteSortByNameActionTagCategorySortCaptionEfter &namnHelpKeywordui_file_panel#sorting_filesHint3   Sortera efter namn|Sortera fjärrpanelen efter namn
ImageIndexShortCutr@  TActionRemoteSortByExtActionTagCategorySortCaption   Efter &filändelseHelpKeywordui_file_panel#sorting_filesHintA   Sortera efter filändelse|Sortera fjärrpanelen efter filändelse
ImageIndex ShortCuts@  TActionRemoteSortBySizeActionTagCategorySortCaptionEfter &storlekHelpKeywordui_file_panel#sorting_filesHint<   Sortera efter storlek|Sortera fjärrpanelen efter filstorlek
ImageIndex#ShortCutu@  TActionRemoteSortByRightsActionTagCategorySortCaption   Efter &filrättigheterHelpKeywordui_file_panel#sorting_filesHintI   Sortera efter filrättigheter|Sortera fjärrpanelen efter filrättigheter
ImageIndex$ShortCutv@  TActionRemoteSortByChangedActionTagCategorySortCaption   Efter senast &ändradHelpKeywordui_file_panel#sorting_filesHintH   Sortera efter senast &ändrad|Sortera fjärrpanelen efter senast ändrad
ImageIndex!ShortCutt@  TActionRemoteSortByOwnerActionTagCategorySortCaption   Efter ä&gareHelpKeywordui_file_panel#sorting_filesHint:   Sortera efter ägare|Sortera fjärrpanelen efter filägare
ImageIndex&ShortCutw@  TActionRemoteSortByGroupActionTagCategorySortCaptionEfter &gruppHelpKeywordui_file_panel#sorting_filesHint8   Sortera efter grupp|Sortera fjärrpanelen efter filgrupp
ImageIndex'ShortCutx@  TActionRemoteSortByTypeActionTagCategorySortCaptionEfter fil&typHelpKeywordui_file_panel#sorting_filesHint7   Sortera efter filtyp|Sortera fjärrkatalog efter filtyp
ImageIndex"  TActionCurrentSortAscendingActionTagCategorySortCaption	Stig&andeHelpKeywordui_file_panel#sorting_filesHintW   Stigande/fallande|Växla sortering mellan stigande och fallande ordning i aktuell panel
ImageIndex%  TActionCurrentSortByNameActionTagCategorySortCaptionEfter &namnHelpKeywordui_file_panel#sorting_filesHint3Sortera efter namn|Sortera aktuell panel efter namn
ImageIndexShortCutr@  TActionCurrentSortByExtActionTagCategorySortCaption   Efter &filändelseHelpKeywordui_file_panel#sorting_filesHintA   Sortera efter filändelse|Sortera aktuell panel efter filändelse
ImageIndex ShortCuts@  TActionCurrentSortBySizeActionTagCategorySortCaptionEfter &storlekHelpKeywordui_file_panel#sorting_filesHint<Sortera efter storlek|Sortera aktuell panel efter filstorlek
ImageIndex#ShortCutu@  TActionCurrentSortByTypeActionTagCategorySortCaptionEfter fil&typHelpKeywordui_file_panel#sorting_filesHintLSortera efter filtyp|Sortera aktuell panel efter filtyp (endast lokal panel)
ImageIndex"  TActionCurrentSortByRightsActionTagCategorySortCaptionEfter &attributHelpKeywordui_file_panel#sorting_filesHintK   Sortera efter attribut|Sortera aktuell panel efter attribut/filrättigheter
ImageIndex$ShortCutv@  TActionCurrentSortByChangedActionTagCategorySortCaption   Efter senast &ändradHelpKeywordui_file_panel#sorting_filesHintH   Sortera efter senast &ändrad|Sortera aktuell panel efter senast ändrad
ImageIndex!ShortCutt@  TActionCurrentSortByOwnerActionTagCategorySortCaption   Efter ä&gareHelpKeywordui_file_panel#sorting_filesHintO   Sortera efter ägare|Sortera aktuell panel efter filägare (endast fjärrpanel)
ImageIndex&ShortCutw@  TActionCurrentSortByGroupActionTagCategorySortCaptionEfter &gruppHelpKeywordui_file_panel#sorting_filesHintM   Sortera efter grupp|Sortera fjärrpanelen efter filgrupp (endast fjärrpanel)
ImageIndex'ShortCutx@  TActionSortColumnAscendingActionTagCategorySortCaptionSortera stig&andeHelpKeywordui_file_panel#sorting_filesHint(Sortera filer stigande efter vald kolumn
ImageIndex)  TActionSortColumnDescendingActionTagCategorySortCaptionSortera fallan&deHelpKeywordui_file_panel#sorting_filesHint(Sortera filer fallande efter vald kolumn
ImageIndex(  TActionHomepageActionTagCategoryHelpCaptionProdukt&hemsidaHint9   Öppnar webbläsaren och går till applikationens hemsida
ImageIndex*  TActionHistoryPageActionTagCategoryHelpCaption&VersionshistorikHintO   Öppnar webbläsaren och går till webbsida med applikationens versionshistorik  TActionSaveCurrentSessionAction2TagCategorySessionCaption&Spara session som webbplats...HelpKeyword&task_connections#saving_opened_sessionHint?Spara session som webbplats|Spara aktuell session som webbplats
ImageIndex+  TActionShowHideRemoteNameColumnActionTagCategoryColumnsCaption&NamnHelpKeywordui_file_panel#selecting_columnsHint5   Visa/dölj namn|Visa/dölj namnkolumn i fjärrpanelen
ImageIndex,  TActionShowHideRemoteExtColumnActionTagCategoryColumnsCaption   &FiländelseHelpKeywordui_file_panel#selecting_columnsHintC   Visa/dölj filändelse|Visa/dölj filändelsekolumn i fjärrpanelen
ImageIndex-  TActionShowHideRemoteSizeColumnActionTagCategoryColumnsCaption&StorlekHelpKeywordui_file_panel#selecting_columnsHint?   Visa/dölj storlek|Visa/dölj filstorlekskolumn i fjärrpanelen
ImageIndex/  TAction!ShowHideRemoteChangedColumnActionTagCategoryColumnsCaption   Se&nast ändradHelpKeywordui_file_panel#selecting_columnsHintJ   Visa/dölj senast ändrad|Visa/dölj senast ändrad-kolumn i fjärrpanelen
ImageIndex0  TAction ShowHideRemoteRightsColumnActionTagCategoryColumnsCaption   Fil&rättigheterHelpKeywordui_file_panel#selecting_columnsHintJ   Visa/dölj filrättigheter|Visa/dölj filrättighetskolumn i fjärrpanelen
ImageIndex1  TActionShowHideRemoteOwnerColumnActionTagCategoryColumnsCaption   &ÄgareHelpKeywordui_file_panel#selecting_columnsHint8   Visa/dölj ägare|Visa/dölj ägarkolumn i fjärrpanelen
ImageIndex2  TActionShowHideRemoteGroupColumnActionTagCategoryColumnsCaption&GruppHelpKeywordui_file_panel#selecting_columnsHint7   Visa/dölj grupp|Visa/dölj gruppkolumn i fjärrpanelen
ImageIndex3  TAction$ShowHideRemoteLinkTargetColumnActionTagCategoryColumnsCaption
   &LänkmålHelpKeywordui_file_panel#selecting_columnsHint@   Visa/dölj länkmål|Visa/dölj länkmålskolumn i fjärrpanelen
ImageIndexR  TActionShowHideRemoteTypeColumnActionTagCategoryColumnsCaptionFil&typHelpKeywordui_file_panel#selecting_columnsHint:   Visa/dölj filtyp|Visa/dölj filtypskolumn i fjärrpanelen
ImageIndex.  TActionShowHideLocalNameColumnActionTagCategoryColumnsCaption&NamnHelpKeywordui_file_panel#selecting_columnsHint:   Visa/dölj namn|Visa/dölj namnkolumn i den lokala panelen
ImageIndex,  TActionShowHideLocalExtColumnActionTagCategoryColumnsCaption   &FiländelseHelpKeywordui_file_panel#selecting_columnsHintH   Visa/dölj filändelse|Visa/dölj filändelsekolumn i den lokala panelen
ImageIndex-  TActionShowHideLocalTypeColumnActionTagCategoryColumnsCaptionFil&typHelpKeywordui_file_panel#selecting_columnsHint?   Visa/dölj filtyp|Visa/dölj filtypskolumn i den lokala panelen
ImageIndex.  TActionShowHideLocalSizeColumnActionTagCategoryColumnsCaption&StorlekHelpKeywordui_file_panel#selecting_columnsHintD   Visa/dölj storlek|Visa/dölj filstorlekskolumn i den lokala panelen
ImageIndex/  TAction ShowHideLocalChangedColumnActionTagCategoryColumnsCaption   Senast &ändradHelpKeywordui_file_panel#selecting_columnsHintO   Visa/dölj senast ändrad|Visa/dölj senast ändrad-kolumn i den lokala panelen
ImageIndex0  TActionShowHideLocalAttrColumnActionTagCategoryColumnsCaption	&AttributHelpKeywordui_file_panel#selecting_columnsHintB   Visa/dölj attribut|Visa/dölj attributkolumn i den lokala panelen
ImageIndex1  TActionCompareDirectoriesActionTagCategoryCommandCaption   &Jämför katalogerHelpKeywordtask_compare_directoriesHintH   Jämför kataloger|Markerar skillnader mellan lokal- och fjärrkatalogen
ImageIndex4ShortCutq   TActionSynchronizeActionTagCategoryCommandCaption!   &Håll fjärrkatalogen uppdateradHelpKeywordtask_keep_up_to_dateHintA   Håll fjärrkatalogen uppdaterad|Håll fjärrkatalogen uppdaterad
ImageIndex5ShortCutU@  TActionForumPageActionTagCategoryHelpCaption&SupportforumHint=   Öppnar webbläsaren och gå till webbsida med supportforumet  TActionLocalAddBookmarkActionTag	CategoryLocal DirectoryCaption   &Lägg till bokmärkenHelpKeywordtask_navigate#bookmarksHintD   Lägg till bokmärken|Lägg till aktuell lokal katalog som bokmärke
ImageIndex6ShortCutB@  TActionRemoteAddBookmarkActionTagCategoryRemote DirectoryCaption   &Lägg till bokmärkenHelpKeywordtask_navigate#bookmarksHintD   Lägg till bokmärken|Lägg till aktuell fjärrkatalog som bokmärke
ImageIndex6ShortCutB@  TActionConsoleActionTagCategoryCommandCaption   Öppna &terminalfönsterHelpKeyword
ui_consoleHint�   Öppna terminalfönster|Öppnar terminalfönster som tillåter körande av godtyckligt extrakommando (med undantag av de som kräver användarinput)
ImageIndex7ShortCutT@  TActionPuttyActionTagCategoryCommandCaption   Öppna session i &PuTTYHelpKeywordintegration_putty#open_puttyHintZ   Öppna session i PuTTY|Starta PuTTY SSH-terminalprogram och öppna aktuell session med den
ImageIndex@ShortCutP@  TActionLocalExploreDirectoryActionTagCategoryLocal DirectoryCaption&Utforska katalogHint+   Öppnar utforskaren i aktuell lokal katalog
ImageIndex8ShortCutE�    TActionCurrentOpenActionTagCategoryFocused OperationCaption   &ÖppnaHelpKeyword	task_editHintQ   Öppna dokument|Öppnar valt dokument med program som filtypen är associerad med
ImageIndex:  TActionSynchronizeBrowsingActionTagCategoryCommand	AutoCheck	Caption   Synkronisera &bläddringHelpKeyword"task_navigate#synchronize_browsingHintJ   Synkronisera bläddring|Synkronisera lokal och fjärrkatalogens bläddring
ImageIndex;ShortCutB�    TActionCurrentAddEditLinkActionTagCategorySelected OperationCaption   Lägg till/redigera &länk...HelpKeyword	task_linkHintZ   Lägg till/redigera länk|Lägger till ny länk/genväg eller redigerar vald länk/genväg
ImageIndex<  TActionCurrentAddEditLinkContextActionTagCategorySelected OperationCaption   Redigera &länk...HelpKeyword	task_linkHint*   Redigera länk|Redigera vald länk/genväg
ImageIndex<  TActionCloseApplicationActionTagCategoryCommandCaption&AvslutaHintG   Avsluta applikation|Avsluta öppnade sessioner och stäng applikationen  TActionOpenedSessionsActionTagCategorySessionCaption   &Öppna sessionerHelpKeyword&task_connections#switching_connectionsHint0   Välj session|Välj öppnad session att aktivera
ImageIndex>  TActionDuplicateSessionActionTagCategorySessionCaption&Dubblera sessionHelpKeywordtask_connectionsHintf   Dubblera session|Öppnar samma session igen (håll nere SHIFT för att öppna den i ett nytt fönster)
ImageIndex[  TActionNewLinkActionTagCategoryCommandCaption	   &Länk...HelpKeyword	task_linkHint"   Skapa länk|Skapa ny länk/genväg
ImageIndex<  TActionCustomCommandsActionTagCategoryCommandCaptionEgna &kommandonHelpKeywordremote_command#custom_commandsHint,   Kör egna kommandon med de markerade filerna  TActionCustomCommandsCustomizeActionTagCategoryCommandCaption&Anpassa...HelpKeywordui_pref_commandsHintAnpassa egna kommandon
ImageIndex  TActionCustomCommandsEnterActionTagCategoryCommandCaption   Lä&gg in...HelpKeyword8remote_command#executing_and_configuring_custom_commandsHint#   Lägg in egna kommandon för ad hoc
ImageIndexZ  TAction CustomCommandsEnterFocusedActionTagCategoryCommandCaption   Lä&gg in...HelpKeyword8remote_command#executing_and_configuring_custom_commandsHint#   Lägg in egna kommandon för ad hoc
ImageIndexZ  TActionCheckForUpdatesActionTagCategoryHelpCaption   Sök efter &uppdateringarHelpKeywordupdatesHint0   Frågar applikationens webbsida om uppdateringar
ImageIndex?  TActionDonatePageActionTagCategoryHelpCaption&DoneraHintG   Öppnar webbläsaren och går till programmets webbsida för donationer  TActionCustomCommandsLastActionTagCategoryCommandCaptionCustomCommandsLastActionHelpKeyword8remote_command#executing_and_configuring_custom_commands  TActionCustomCommandsLastFocusedActionTagCategoryCommandCaptionCustomCommandsLastFocusedActionHelpKeyword8remote_command#executing_and_configuring_custom_commands  TActionFileSystemInfoActionTagCategoryCommandCaption&Server/protokollinformationHelpKeyword	ui_fsinfoHint Visa server/protokollinformation
ImageIndex  TActionClearCachesActionTagCategoryCommandCaption&Rensa cacheHelpKeyworddirectory_cacheHint1   Rensa cache för kataloglistning och katalogbyten  TActionFullSynchronizeActionTagCategoryCommandCaption&Synkronisera...HelpKeywordtask_synchronize_fullHint,   Synkronisera lokal katalog med fjärrkatalog
ImageIndexBShortCutS@  TActionRemoteMoveToFocusedActionTagCategoryRemote Focused OperationCaption&Flytta till...HelpKeyword'task_move_duplicate#moving_remote_filesHint0   Flytta|Flytta markerade filer till fjärrkatalog
ImageIndexd  TActionShowHiddenFilesActionTagCategoryViewCaption   Visa/dölj &dolda filerHelpKeywordui_file_panel#special_filesHint)   Växla visning av dolda filer i panel(er)ShortCutH�    TActionFormatSizeBytesActionTagCategoryViewCaptionKorta &filstorlekarHelpKeywordui_file_panel#short_formatHint-Visa filstorlekar i kort format (kB, MB, etc)  TActionLocalPathToClipboardActionTagCategoryLocal DirectoryCaption   Kopiera s&ökväg till urklippHelpKeyword#filenames#current_working_directoryHint+   Kopiera aktuell lokal sökväg till urklipp  TActionRemotePathToClipboardActionTagCategoryRemote DirectoryCaption   Kopiera s&ökväg till urklippHelpKeyword#filenames#current_working_directoryHint+   Kopiera aktuell fjärrsökväg till urklipp  TActionFileListToCommandLineActionTagCategorySelected OperationCaptionIn&foga till kommandoradHelpKeywordfilenames#command_lineHint/Infoga markerade filers namn till kommandoradenShortCut@  TActionFileListToClipboardActionTagCategorySelected OperationCaption&Kopiera till urklippHelpKeywordfilenames#file_nameHint*Kopiera markerade filers namn till urklippShortCutC`  TActionFullFileListToClipboardActionTagCategorySelected OperationCaption,   Kopiera till urklipp (inklusive s&ökvägar)HelpKeywordfilenames#file_nameHint=   Kopiera markerade filers namn inklusive sökväg till urklippShortCutC�    TActionQueueGoToActionTagCategoryQueueCaption	   &Gå tillHelpKeywordui_queue#managing_the_queueHint   Gå till överföringskölistan
ImageIndexJShortCutQ@  TActionQueueItemUpActionTagCategoryQueueCaptionFlytta &uppHelpKeywordui_queue#managing_the_queueHint2   Flytta upp vald köpost för att utföras tidigare
ImageIndexH  TActionQueueItemDownActionTagCategoryQueueCaptionFlytta &nerHelpKeywordui_queue#managing_the_queueHint0   Flytta ner vald köpost för att utföras senare
ImageIndexI  TActionQueueToggleShowActionTagCategoryQueueCaption   &KöHint   Visa/dölj kölista
ImageIndexJ  TActionQueueShowActionTagCategoryQueueCaptionVi&saHelpKeywordui_queueHint   Visa kölista  TActionQueueHideWhenEmptyActionTagCategoryQueueCaption   Dölj ifall &tomHelpKeywordui_queueHint    Dölj kölistan när den är tom  TActionQueueHideActionTagCategoryQueueCaption   &DöljHelpKeywordui_queueHint   Dölj kölista  TActionQueueToolbarActionTagCategoryQueueCaption   &VerktygsfältHint@   Dölj/visa verktygsfältet för kölistan (på kölistans panel)  TActionQueuePreferencesActionTagCategoryQueueCaptionA&npassa...HelpKeywordui_pref_backgroundHint   Anpassa kölista
ImageIndex  TActionPasteActionTagCategoryCommandCaptionK&listra inHelpKeyword task_upload#using_copy_amp:pasteHintA   Klistra in filer från urklipp till aktuell katalog i aktiv panel
ImageIndexKShortCutV@  TActionNewFileActionTagCategoryCommandCaption&Fil...HelpKeyword	task_editHint1   Skapa fil|Skapar ny fil och öppnas den i editorn
ImageIndexM  TActionEditorListCustomizeActionTagCategoryCommandCaption&Konfigurera...HelpKeywordui_pref_editorHint   Skräddarsy editorer
ImageIndex  TActionRemoteCopyToFocusedActionTagCategoryRemote Focused OperationCaption&Dubblera...HelpKeyword,task_move_duplicate#duplicating_remote_filesHint3   Dubblera|Dubbleras valda filer till fjärrkatalogen
ImageIndexN  TActionRemoteCopyToActionTagCategoryRemote Selected OperationCaption&Dubblera...HelpKeyword,task_move_duplicate#duplicating_remote_filesHint2   Dubblera|Dubblera valda filer till fjärrkatalogen
ImageIndexN  TActionUrlToClipboardActionTagCategorySelected OperationCaptionKopiera &URL till urklippHelpKeywordfilenames#file_urlHint*Kopiera URL'er av valda filer till urklipp  TActionTableOfContentsActionTagCategoryHelpCaption
   I&nnehållHintI   Öppnar webbläsare och går till dokumentationens innehållsförteckning
ImageIndexOShortCutp  TActionFileListFromClipboardActionTagCategorySelected OperationCaption&Transfer Files in ClipboardHint+Transfer files whose names are in clipboard  TActionLocalCopyActionTag	CategoryLocal Selected OperationCaption   &Överför...HelpKeywordtask_uploadHint   Överför|Överför valda filer
ImageIndexX  TActionCurrentDeleteAlternativeActionTagCategorySelected OperationCaption&Ta bortHelpKeywordtask_deleteHintTa bort|Ta bort valda filer
ImageIndex  TActionCurrentEditAlternativeActionTagCategorySelected OperationCaption&Redigera (alternativ)HelpKeyword	task_editHint@Redigera (alternativ)|Redigera valda filer med alternativ editor  TActionCurrentEditWithActionTagCategorySelected OperationCaptionRedigera &med...HelpKeyword	task_editHint9Redigera med|Redigera valda filer med editorn som ni valt  TActionDownloadPageActionTagCategoryHelpCaption
Ladda &nerHintA   Öppnar webbläsare och går till applikationens nerladdningssida  TActionUpdatesPreferencesActionTagCategoryHelpCaptionKonfi&gurera...HelpKeywordui_pref_updatesHintC   Konfigurera automatisk kontroll av uppdateringar för applikationen
ImageIndex  TActionShowUpdatesActionTagCategoryHelpCaption&Visa uppdateringarHelpKeywordupdatesHint�   Visa information om applikationens uppdateringar|Visa information om applikationens uppdateringar (förfrågar applikationens hemsida om informationen inte är tillgänglig vid tidpunkten)
ImageIndexQ  TActionPresetsPreferencesActionTagCategoryViewCaption&Konfigurera...HelpKeywordui_pref_presetsHint2   Konfigurera förinställningar för överföringar
ImageIndex  TActionLockToolbarsActionTagCategoryViewCaption   &Lås verktygsfältHelpKeywordui_toolbarsHint3   Hindra flyttning och dockning av alla verktygsfält  TActionSelectiveToolbarTextActionTagCategoryViewCaption&Visa valbara textetiketterHelpKeywordui_toolbarsHintD   Visa textetiketter på utvalda viktiga kommandon på verktygsfältet  TActionCustomCommandsBandActionTagCategoryViewCaptionEgna ko&mmandoknapparHelpKeywordui_toolbarsHint,   Dölj/visa verktygsfält för egna kommandon  TActionColorMenuActionTagCategoryViewCaption   F&ärgHelpKeywordtask_connections#session_colorHint    Ändra färg på aktuell session  TActionAutoReadDirectoryAfterOpActionTagCategoryViewCaptionLadda auto&matisk om katalogHint=   Ändra automatisk omladdning av fjärrkatalog efter operationShortCutR�    TActionQueueItemPauseActionTagCategoryQueueCaption&PausaHelpKeywordui_queue#managing_the_queueHint   Pausa vald köpost
ImageIndexS  TActionQueueItemResumeActionTagCategoryQueueCaption   &ÅterupptaHelpKeywordui_queue#managing_the_queueHint   Återuppta vald pausad köpost
ImageIndexF  TActionQueuePauseAllActionTagCategoryQueueCaption&Pausa allaHelpKeywordui_queue#managing_the_queueHint   Pausa alla köposter som körs
ImageIndexT  TActionQueueResumeAllActionTagCategoryQueueCaption   &Återuppta allaHelpKeywordui_queue#managing_the_queueHint!   Återuppta alla pausade köposter
ImageIndexU  TActionQueueDeleteAllDoneActionTagCategoryQueueCaption   Ta bort alla &slutfördaHelpKeywordui_queue#managing_the_queueHint!   Ta bort alla slutförda köposter
ImageIndexc  TActionQueueEnableActionTagCategoryQueueCaption   &ProcessköHelpKeywordui_queue#managing_the_queueHints   Aktivera köbehandling|Aktivera köbehandling (väntande köposter startar inte, när köbehandling är inaktiverad
ImageIndex`ShortCutQ`  TActionQueueDisconnectOnceEmptyActionTagCategoryQueueCaption   &Koppla ifrånHelpKeywordui_queueHint'   Koppla ifrån session när kön är tom
ImageIndexW  TActionRestoreSelectionActionTagCategory	SelectionCaption   &Återställ markeringHelpKeywordui_file_panel#selecting_filesHint"   Återställ föregående markering
ImageIndexV  TActionLocalSelectActionTagCategory	SelectionCaption&Markera filerHelpKeyword	ui_selectHint'Markera|Markera lokala filer efter mask
ImageIndex  TActionLocalUnselectActionTagCategory	SelectionCaptionA&vmarkera filerHelpKeyword	ui_selectHint+Avmarkera|Avmarkera lokala filer efter mask
ImageIndex  TActionLocalSelectAllActionTagCategory	SelectionCaptionM&arkera allaHelpKeywordui_file_panel#selecting_filesHintMarkera alla lokala filer
ImageIndex  TActionCurrentEditFocusedActionTagCategoryFocused OperationCaption	&RedigeraHelpKeyword	task_editHintRedigera|Redigera valda filer
ImageIndex9  TActionNewDirActionTagCategoryCommandCaptionKatalo&g...HelpKeywordtask_create_directoryHintSkapa katalog|Skapa ny katalog
ImageIndex  TActionQueueShutDownOnceEmptyActionTagCategoryQueueCaption   &Sträng av datornHelpKeywordui_queueHint#   Sträng av datorn när kön är tom
ImageIndex]  TActionQueueIdleOnceEmptyActionTagCategoryQueueCaption   &Förbli idleChecked	HelpKeywordui_queueHint   Förbli idle när kön är tom
ImageIndex^  TActionQueueCycleOnceEmptyActionTagCategoryQueueCaption   &Tom köHelpKeywordui_queueHint1   Ändra åtgärd som ska utföras då kön är tom
ImageIndex^  TTBEditActionQueueItemSpeedActionTagCategoryQueueHelpKeywordui_queue#managing_the_queueHint)   Ändra hastighetsgräns för vald köpostEditCaption
&Hastighet  TActionLocalFilterActionTag	CategoryLocal DirectoryCaption&Filtrera...HelpKeywordui_file_panel#filterHintFiltrera|Filtrera visade filer
ImageIndex\  TActionRemoteFilterActionTagCategoryRemote DirectoryCaption
&Filter...HelpKeywordui_file_panel#filterHintFilter|Filtrera visade filer
ImageIndex\  TActionRemoteFindFilesActionTagCategoryRemote DirectoryCaption   Sö&k filer..HelpKeyword	task_findHint#   Sök filer|Sök filer och kataloger
ImageIndex_  TActionCurrentEditInternalActionTagCategorySelected OperationCaption&Intern editorHelpKeyword	task_editHint8Redigera (intern)|Redigera valda filer med intern editor  TActionSaveWorkspaceActionTagCategorySessionCaptionSpara arbets&yta...HelpKeyword	workspaceHintSpara arbetsyta|Spara arbetsyta
ImageIndexf  TActionLocalRenameActionTagCategoryLocal Selected OperationCaption	&Byt namnHelpKeywordtask_renameHint$   Byt namn|Byt namn på vald lokal fil
ImageIndex  TActionLocalEditActionTagCategoryLocal Selected OperationCaption	&RedigeraHelpKeyword	task_editHint$Redigera|Redigera valda lokala filer
ImageIndex9  TActionLocalMoveActionTag	CategoryLocal Selected OperationCaption   Överför och ta &bort...HelpKeywordtask_uploadHint]   Överför och ta bort|Överför valda lokala filer till fjärrkatalogen och tar bort original
ImageIndexb  TActionLocalCreateDirActionTagCategoryLocal Selected OperationCaptionS&kapa katalog...HelpKeywordtask_create_directoryHint$Skapa katalog|Skapa ny lokal katalog
ImageIndex  TActionLocalDeleteActionTagCategoryLocal Selected OperationCaption&Ta bortHelpKeywordtask_deleteHint"Ta bort|Ta bort valda lokala filer
ImageIndex  TActionLocalPropertiesActionTagCategoryLocal Selected OperationCaption&EgenskaperHelpKeywordtask_propertiesHint9   Egenskaper|Visa/ändra egenskaper för valda lokala filer
ImageIndex  TActionLocalAddEditLinkActionTagCategoryLocal Selected OperationCaption   Lägg till/redigera &länk...HelpKeyword	task_linkHint\   Lägg till/redigera genväg|Lägg till en ny lokal genväg eller redigera vald lokal genväg
ImageIndex<  TActionRemoteRenameActionTagCategoryRemote Selected OperationCaption	&Byt namnHelpKeywordtask_renameHint$   Byt namn|Byt namn på vald fjärrfil
ImageIndex  TActionRemoteEditActionTagCategoryRemote Selected OperationCaption	&RedigeraHelpKeyword	task_editHint#   Redigera|Redigera valda fjärrfiler
ImageIndex9  TActionRemoteMoveActionTagCategoryRemote Selected OperationCaptionLadda ner och &ta bortHelpKeywordtask_downloadHintY   Ladda ner och ta bort|Ladda ner valda fjärrfiler till lokal katalog och ta bort original
ImageIndexa  TActionRemoteCreateDirActionTagCategoryRemote Selected OperationCaptionS&kapa katalog...HelpKeywordtask_create_directoryHint$   Skapa katalog|Skapa ny fjärrkatalog
ImageIndex  TActionRemoteDeleteActionTagCategoryRemote Selected OperationCaption&Ta bortHelpKeywordtask_deleteHint!   Ta bort|Ta bort valda fjärrfiler
ImageIndex  TActionRemotePropertiesActionTagCategoryRemote Selected OperationCaption&EgenskaperHelpKeywordtask_propertiesHintZ   Egenskaper|Visa/ändra rättigheter, ägarskap och andra egenskaper för valda fjärrfiler
ImageIndex  TActionRemoteAddEditLinkActionTagCategoryRemote Selected OperationCaption   Lägg till/redigera &länk...HelpKeyword	task_linkHintQ   Lägg till/ändra länk|Lägg till ny fjärrlänk eller redigera vald fjärrlänk
ImageIndex<  TActionRemoteSelectActionTagCategory	SelectionCaption&Markera filerHelpKeyword	ui_selectHint&   Markera|Markera fjärrfiler efter mask
ImageIndex  TActionRemoteUnselectActionTagCategory	SelectionCaptionA&vmarkera filerHelpKeyword	ui_selectHint*   Avmarkera|Avmarkera fjärrfiler efter mask
ImageIndex  TActionRemoteSelectAllActionTagCategory	SelectionCaptionM&arkera allaHelpKeywordui_file_panel#selecting_filesHint   Markera alla fjärrfiler
ImageIndex  TActionLocalMoveFocusedActionTagCategoryLocal Focused OperationCaption   Överför och &ta bort...HelpKeywordtask_uploadHintZ   Överför och ta bort|Överför valda lokala filer till fjärrkatalog och ta bort original
ImageIndexb  TActionCurrentSystemMenuFocusedActionTagCategoryFocused OperationCaption&SystemmenyHintn   Visa filsystemets snabbmeny (i egenskaper kan du välja att visa den som standard istället för inbyggd meny)   TTBXPopupMenuExplorerBarPopupImagesGlyphsModule.ExplorerImagesLeft� TopP TTBXItemAddress2ActionExplorerAddressBandAction  TTBXItemStandardButtons1ActionExplorerToolbarBandAction  TTBXItemSelectionButtons1ActionExplorerSelectionBandAction  TTBXItemSessionButtons2ActionExplorerSessionBandAction  TTBXItemPreferencesButtons1ActionExplorerPreferencesBandAction  TTBXItemSortButtons3ActionExplorerSortBandAction  TTBXItemTBXItem3ActionExplorerUpdatesBandAction  TTBXItemTBXItem4ActionExplorerTransferBandAction  TTBXItem	TBXItem16Action ExplorerCustomCommandsBandAction  TTBXItemTBXItem7ActionLockToolbarsAction  TTBXItem	TBXItem48ActionSelectiveToolbarTextAction  TTBXSeparatorItemN5  TTBXItemSessionsTabsAction2ActionSessionsTabsAction  TTBXItem
StatusBar2ActionStatusBarAction  TTBXSeparatorItemN72  TTBXSubmenuItemQueue7Caption   &KöHelpKeywordui_queueHint   Konfigurera kölista TTBXItemShow6ActionQueueShowAction	RadioItem	  TTBXItemHidewhenEmpty6ActionQueueHideWhenEmptyAction	RadioItem	  TTBXItemHide5ActionQueueHideAction	RadioItem	  TTBXSeparatorItemN71  TTBXItemToolbar5ActionQueueToolbarAction  TTBXSeparatorItemN70  TTBXItem
Customize5ActionQueuePreferencesAction   TTBXItemTree4ActionRemoteTreeAction   TTimerSessionIdleTimerEnabledInterval�OnTimerSessionIdleTimerTimerLeft TopP  TTBXPopupMenuCommanderBarPopupImagesGlyphsModule.ExplorerImagesLeft�Top TTBXItemCommandsButtons2ActionCommanderCommandsBandAction  TTBXItemSessionButtons5ActionCommanderSessionBandAction  TTBXItemPreferencesButtons4ActionCommanderPreferencesBandAction  TTBXItemSortButtons2ActionCommanderSortBandAction  TTBXItemTBXItem2ActionCommanderUpdatesBandAction  TTBXItemTBXItem5ActionCommanderTransferBandAction  TTBXItem	TBXItem15Action!CommanderCustomCommandsBandAction  TTBXItemTBXItem6ActionLockToolbarsAction  TTBXItem	TBXItem46ActionSelectiveToolbarTextAction  TTBXSeparatorItemN26  TTBXItemSessionsTabsAction1ActionSessionsTabsAction  TTBXItemCommandLine2ActionCommandLinePanelAction  TTBXItemCommandsToolbar1ActionToolBar2Action  TTBXItem
StatusBar8ActionStatusBarAction  TTBXSeparatorItemN27  TTBXSubmenuItemLocalPanel1Caption&Lokal panelHelpKeywordui_file_panelHint#   Ändra den lokala panelens utseende TTBXItemHistoryButtons3ActionCommanderLocalHistoryBandAction  TTBXItemNavigationButtons3Action"CommanderLocalNavigationBandAction  TTBXItem	TBXItem40ActionCommanderLocalFileBandAction  TTBXItem	TBXItem43Action!CommanderLocalSelectionBandAction  TTBXSeparatorItemN23  TTBXItemTree7ActionLocalTreeAction  TTBXSeparatorItemN77  TTBXItem
StatusBar6ActionLocalStatusBarAction   TTBXSubmenuItemRemotePanel2Caption   &FjärrpanelHelpKeywordui_file_panelHint   Ändra fjärrpanelens utseende TTBXItemHistoryButtons4Action CommanderRemoteHistoryBandAction  TTBXItemNavigationButtons4Action#CommanderRemoteNavigationBandAction  TTBXItem	TBXItem41ActionCommanderRemoteFileBandAction  TTBXItem	TBXItem42Action"CommanderRemoteSelectionBandAction  TTBXSeparatorItemN25  TTBXItemTree8ActionRemoteTreeAction  TTBXSeparatorItemN78  TTBXItem
StatusBar7ActionRemoteStatusBarAction   TTBXSubmenuItemOptions1Caption   &KöHelpKeywordui_queueHint   Konfigurera kölista TTBXItemShow5ActionQueueShowAction	RadioItem	  TTBXItemHidewhenEmpty5ActionQueueHideWhenEmptyAction	RadioItem	  TTBXItemHide4ActionQueueHideAction	RadioItem	  TTBXSeparatorItemN69  TTBXItemToolbar4ActionQueueToolbarAction  TTBXSeparatorItemN68  TTBXItem
Customize4ActionQueuePreferencesAction    TTBXPopupMenuRemotePanelPopupImagesGlyphsModule.ExplorerImagesLeft8Top TTBXItem	TBXItem32ActionRemoteRefreshAction  TTBXItem	TBXItem30ActionRemoteAddBookmarkAction  TTBXItemCopyPathtoClipboard1ActionRemotePathToClipboardAction  TTBXItemOpenDirectoryBookmark1ActionRemoteOpenDirAction  TTBXItem	TBXItem26ActionRemoteFilterAction  TTBXSeparatorItemN51  TTBXItemHistoryButtons5Action CommanderRemoteHistoryBandAction  TTBXItemNavigationButtons5Action#CommanderRemoteNavigationBandAction  TTBXItem	TBXItem14ActionCommanderRemoteFileBandAction  TTBXItem	TBXItem45Action"CommanderRemoteSelectionBandAction  TTBXItem	TBXItem37ActionLockToolbarsAction  TTBXItem	TBXItem49ActionSelectiveToolbarTextAction  TTBXSeparatorItemN28  TTBXItemTree5ActionRemoteTreeAction  TTBXSeparatorItemN75  TTBXItem
StatusBar9ActionRemoteStatusBarAction   TTBXPopupMenuLocalPanelPopupImagesGlyphsModule.ExplorerImagesLeft8TopP TTBXItem	TBXItem34ActionLocalRefreshAction  TTBXItem	TBXItem31ActionLocalAddBookmarkAction  TTBXItemCopyPathtoClipboard2ActionLocalPathToClipboardAction  TTBXItemOpenDirectoryBookmark2ActionLocalOpenDirAction  TTBXItem	TBXItem27ActionLocalFilterAction  TTBXSeparatorItemN52  TTBXItemHistoryButtons6ActionCommanderLocalHistoryBandAction  TTBXItemNavigationButtons6Action"CommanderLocalNavigationBandAction  TTBXItem	TBXItem39ActionCommanderLocalFileBandAction  TTBXItem	TBXItem44Action!CommanderLocalSelectionBandAction  TTBXItem	TBXItem38ActionLockToolbarsAction  TTBXItem	TBXItem47ActionSelectiveToolbarTextAction  TTBXSeparatorItemN29  TTBXItemTree6ActionLocalTreeAction  TTBXSeparatorItemN76  TTBXItemStatusBar10ActionLocalStatusBarAction   TTBXPopupMenuLocalDirViewColumnPopupImagesGlyphsModule.ExplorerImagesLeft� TopX TTBXItemSortAscending1ActionSortColumnAscendingAction  TTBXItemSortDescending1ActionSortColumnDescendingAction  TTBXItemLocalSortByExtColumnPopupItemActionLocalSortByExtAction  TTBXItemLocalFormatSizeBytesPopupItemActionFormatSizeBytesAction  TTBXItemHidecolumn1ActionHideColumnAction  TTBXSeparatorItemN37  TTBXSubmenuItemShowcolumns3CaptionVisa &kolumnerHelpKeywordui_file_panel#selecting_columnsHint&   Välj kolumner som ska visas i panelen TTBXItemName3ActionShowHideLocalNameColumnAction  TTBXItemSize3ActionShowHideLocalSizeColumnAction  TTBXItemType2ActionShowHideLocalTypeColumnAction  TTBXItemModification3Action ShowHideLocalChangedColumnAction  TTBXItemAttributes3ActionShowHideLocalAttrColumnAction    TTBXPopupMenuRemoteDirViewColumnPopupImagesGlyphsModule.ExplorerImagesLeft�TopX TTBXItem	MenuItem1ActionSortColumnAscendingAction	RadioItem	  TTBXItem	MenuItem2ActionSortColumnDescendingAction	RadioItem	  TTBXItemRemoteSortByExtColumnPopupItemActionRemoteSortByExtAction  TTBXItemRemoteFormatSizeBytesPopupItemActionFormatSizeBytesAction  TTBXItemHidecolumn2ActionHideColumnAction  TTBXSeparatorItemN38  TTBXSubmenuItemShowcolumns4CaptionVisa &kolumnerHelpKeywordui_file_panel#selecting_columnsHint&   Välj kolumner som ska visas i panelen TTBXItemName4ActionShowHideRemoteNameColumnAction  TTBXItemSize4ActionShowHideRemoteSizeColumnAction  TTBXItemTBXItem8ActionShowHideRemoteTypeColumnAction  TTBXItemModification4Action!ShowHideRemoteChangedColumnAction  TTBXItemPermissions1Action ShowHideRemoteRightsColumnAction  TTBXItemOwner2ActionShowHideRemoteOwnerColumnAction  TTBXItemGroup2ActionShowHideRemoteGroupColumnAction  TTBXItemTBXItem1Action$ShowHideRemoteLinkTargetColumnAction    TTBXPopupMenu
QueuePopupImagesGlyphsModule.ExplorerImagesOnPopupQueuePopupPopupLeft�Top�  TTBXItem
ShowQuery1ActionQueueItemQueryAction  TTBXItem
ShowError1ActionQueueItemErrorAction  TTBXItemShowPrompt1ActionQueueItemPromptAction  TTBXSeparatorItemN53  TTBXItemExecuteNow1ActionQueueItemExecuteAction  TTBXItemTBXItem9ActionQueueItemPauseAction  TTBXItem	TBXItem10ActionQueueItemResumeAction  TTBXItemDelete4ActionQueueItemDeleteAction  TTBXComboBoxItemQueuePopupSpeedComboBoxItemActionQueueItemSpeedAction  TTBXSeparatorItemN54  TTBXItemMoveUp1ActionQueueItemUpAction  TTBXItem	MoveDown1ActionQueueItemDownAction  TTBXSeparatorItemN67  TTBXItemQueueEnableItemActionQueueEnableAction  TTBXSubmenuItemTBXSubmenuItem1Caption&AllaHelpKeywordui_queue#managing_the_queueHint&   Administrationskommandon för kömassa TTBXItem	TBXItem11ActionQueuePauseAllAction  TTBXItem	TBXItem12ActionQueueResumeAllAction  TTBXSeparatorItemTBXSeparatorItem5  TTBXItem	TBXItem51ActionQueueDeleteAllDoneAction   TTBXSubmenuItemTBXSubmenuItem3ActionQueueCycleOnceEmptyActionDropdownCombo	 TTBXItem	TBXItem28ActionQueueIdleOnceEmptyAction	RadioItem	  TTBXItem	TBXItem13ActionQueueDisconnectOnceEmptyAction	RadioItem	  TTBXItem	TBXItem29ActionQueueShutDownOnceEmptyAction	RadioItem	   TTBXSubmenuItemQueue2Caption&AlternativHelpKeywordui_queueHint   Konfigurera kölista TTBXItemShow4ActionQueueShowAction	RadioItem	  TTBXItemHidewhenEmpty4ActionQueueHideWhenEmptyAction	RadioItem	  TTBXItemHide3ActionQueueHideAction	RadioItem	  TTBXSeparatorItemN66  TTBXItemToolbar3ActionQueueToolbarAction  TTBXSeparatorItemN65  TTBXItem
Customize3ActionQueuePreferencesAction    TTBXPopupMenuRemoteDirViewPopup	AutoPopupImagesGlyphsModule.ExplorerImagesLefthTop� TTBXSubmenuItemGoTo4Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItemOpenDirectoryBookmark3ActionRemoteOpenDirAction  TTBXSeparatorItemN81  TTBXItemParentDirectory4ActionRemoteParentDirAction  TTBXItemRootDirectory4ActionRemoteRootDirAction  TTBXItemHomeDirectory4ActionRemoteHomeDirAction  TTBXSeparatorItemN80  TTBXItemBack4ActionRemoteBackAction  TTBXItemForward4ActionRemoteForwardAction   TTBXItemRefresh4ActionRemoteRefreshAction  TTBXItemAddToBookmarks4ActionRemoteAddBookmarkAction  TTBXItem	TBXItem35ActionRemoteFilterAction  TTBXItemCopyPathtoClipboard6ActionRemotePathToClipboardAction  TTBXSeparatorItemN79  TTBXSubmenuItemTBXSubmenuItem26Caption&NyHelpKeyword
task_indexHintSkapa objekt|Skapa nytt objekt TTBXItem
TBXItem135ActionNewFileAction  TTBXItem
TBXItem136ActionNewDirAction  TTBXItem
TBXItem209ActionNewLinkAction    TTBXPopupMenuLocalDirViewPopup	AutoPopupImagesGlyphsModule.ExplorerImagesLeft�Top� TTBXSubmenuItemGoTo5Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItemOpenDirectoryBookmark4ActionLocalOpenDirAction  TTBXItemExploreDirectory2ActionLocalExploreDirectoryAction  TTBXSeparatorItemN84  TTBXItemParentDirectory5ActionLocalParentDirAction  TTBXItemRootDirectory5ActionLocalRootDirAction  TTBXItemHomeDirectory5ActionLocalHomeDirAction  TTBXSeparatorItemN83  TTBXItemBack5ActionLocalBackAction  TTBXItemForward5ActionLocalForwardAction   TTBXItemRefresh5ActionLocalRefreshAction  TTBXItem	TBXItem36ActionLocalFilterAction  TTBXItemAddToBookmarks5ActionLocalAddBookmarkAction  TTBXItemCopyPathtoClipboard7ActionLocalPathToClipboardAction  TTBXSeparatorItemN82  TTBXItemCreateDirectory4ActionCurrentCreateDirAction   TTBXPopupMenuRemoteAddressPopupImagesGlyphsModule.ExplorerImagesLeft� Top� TTBXItem	TBXItem33ActionRemoteRefreshAction  TTBXItem	TBXItem24ActionRemoteAddBookmarkAction  TTBXItem	TBXItem25ActionRemotePathToClipboardAction  TTBXSeparatorItemTBXSeparatorItem1  TTBXItem	TBXItem17ActionRemoteOpenDirAction  TTBXSubmenuItemTBXSubmenuItem2Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItem	TBXItem18ActionRemoteParentDirAction  TTBXItem	TBXItem19ActionRemoteRootDirAction  TTBXItem	TBXItem20ActionRemoteHomeDirAction  TTBXSeparatorItemTBXSeparatorItem2  TTBXItem	TBXItem21ActionRemoteBackAction  TTBXItem	TBXItem22ActionRemoteForwardAction    TTBXPopupMenuSessionsPopupImagesGlyphsModule.ExplorerImagesLeft�Top�  TTBXItem
TBXItem124ActionCloseSessionAction  TTBXItem
TBXItem219ActionDuplicateSessionAction  TTBXItem
TBXItem125ActionSaveCurrentSessionAction2  TTBXSeparatorItemTBXSeparatorItem34  TTBXItem
TBXItem123ActionNewSessionAction  TTBXSubmenuItemTBXSubmenuItem23ActionSavedSessionsAction2OptionstboDropdownArrow   TTBXSeparatorItemTBXSeparatorItem52  TTBXColorItemColorMenuItemActionColorMenuActionColorclNone  TTBXSeparatorItemTBXSeparatorItem35  TTBXItemSessionsTabsAction4ActionSessionsTabsAction   TShellResourcesShellResourcesLeft0Top�  TTBXPopupMenuLocalFilePopupImagesGlyphsModule.ExplorerImagesLeftTopP TTBXItemLocalOpenMenuItemActionCurrentOpenAction  TTBXItemLocalEditMenuItemActionCurrentEditFocusedAction  TTBXItemLocalCopyMenuItemActionLocalCopyFocusedAction  TTBXItem	TBXItem54ActionLocalMoveFocusedAction  TTBXItem	TBXItem57ActionCurrentDeleteFocusedAction  TTBXItem	TBXItem58ActionCurrentRenameAction  TTBXSeparatorItemTBXSeparatorItem3  TTBXSubmenuItemTBXSubmenuItem4ActionCustomCommandsAction TTBXItem    TTBXSubmenuItemTBXSubmenuItem5Caption&FilnamnHelpKeyword	filenamesHint$   Operationer med namn på valda filer TTBXItem	TBXItem59ActionFileListToCommandLineAction  TTBXItem	TBXItem60ActionFileListToClipboardAction  TTBXItem	TBXItem61ActionFullFileListToClipboardAction  TTBXItem	TBXItem62ActionUrlToClipboardAction   TTBXSeparatorItemTBXSeparatorItem4  TTBXItem	TBXItem63ActionCurrentPropertiesFocusedAction  TTBXItem	TBXItem50ActionCurrentSystemMenuFocusedAction       TPF0TOpenDirectoryDialogOpenDirectoryDialogLeft�Top� HelpType	htKeywordHelpKeyword
ui_opendirBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionOpen directoryClientHeightNClientWidth�Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnShowFormShow
DesignSize�N PixelsPerInch`
TextHeight TLabel	EditLabelLeft.TopWidthLHeightCaption   &Öppna katalog:  TImageImageLeftTopWidth Height AutoSize	Picture.Data
*  	TPngImage�PNG

   IHDR           szz�   	pHYs  �  ��o�d  �IDATx��{L[Uǿ����e�.��X��P������l��F�4`��b��l#օ�(�m�_��h�7a5Ƃc�=�M�ɻ��aK�V�����ʥ��1����9���9����~���a4X#����#�=�j���]�3��J��M��� ���wLc��}�ɂ��ާJ��aY� �H�DkfS���Oh�' Q����8�P p��ÿ#nLx����
�^o��\7���ژ�'�Ts�t���
+Xe�����cN�ɉ۸��mR�������.��2>�}��(�O2h�����J�I�D�>��*NC��PA���vv׀�j�PO*+����&ĕV��g<רJ�Y�{������pc�Ht��8��z<k�Z��Sq�ĝە�t�Kj��J_<d,<,+?`�C������;/p<k�!����{��Q�Q��dDr:+;�h��,�)i�Ԋg_��q}�:^�Zz�i���eSX�j<�L��	~��˂�\�L���R7���������K-�w�F j�:�ʶfoڲa������%c� ����O��ܜ��+^\�Ͷ�( r�:o�5)ioX;q����}�l�͉G�eX4٬� �_2�
���hpN,�#"["x^�* ���S�sJ
_��ٹö�#ck�2��)L��� B��y�]��w��N�p�������$ ��C�x���ض�-`����G"��qԜϬ��yF&���y�:�/�Y `�&����`0e���)�T��X���1t�:NP�j	@IA� ��G����zH(�\�o��ˏ�NH ��׺���:��e�:u?�Pt?���3���+���H �41�ڣ��7���Nb���(�
-�(�8�mo(>�hJ-�i	@f�1���ʃ��5��"|,�CmD�tk�sC���f�� RX����,����y�;dQ��m��ƿ.�q���aa,ޅ�i*zܐ�ߜ��N�� ��}�CG�G�y���ďR�'�!�b�I�g�Z�=p��v��8~�`�ў�Jp�,��J�ZP#1����`��ː;
`���� N����Ő����� "~��"l�|N���y]	�f�	����Sr�hc�P*B"ZX�D$�sӅ?���w�Y k��d�=OB��b H�r�R���7(~@���T��:]jL�-��p}8�����Q���(��ڴa�k����a���V��j���FT��5�    IEND�B`�  TIEComboBoxLocalDirectoryEditLeft.TopWidthHeightAnchorsakLeftakTopakRight TabOrderTextLocalDirectoryEditOnChangeDirectoryEditChange  TIEComboBoxRemoteDirectoryEditLeft.TopWidth_HeightAnchorsakLeftakTopakRight 	MaxLength�TabOrder TextRemoteDirectoryEditOnChangeDirectoryEditChange  TButtonOKBtnLeft� Top,WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft� Top,WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TPageControlPageControlLeftTop8Width�Height� 
ActivePageSessionBookmarksSheetAnchorsakLeftakTopakRightakBottom TabOrderOnChangePageControlChange 	TTabSheetSessionBookmarksSheetTagCaption   Sessionsbokmärken
DesignSizez�   TListBoxSessionBookmarksListTagLeft
Top	WidthHeight� AnchorsakLeftakTopakRightakBottom DragModedmAutomatic
ItemHeightTabOrder OnClickBookmarksListClick
OnDblClickBookmarksListDblClick
OnDragDropBookmarksListDragDrop
OnDragOverBookmarksListDragOver	OnEndDragBookmarksListEndDrag	OnKeyDownBookmarksListKeyDownOnStartDragBookmarksListStartDrag  TButtonAddSessionBookmarkButtonTagLeftTop	WidthSHeightAnchorsakTopakRight Caption   &Lägg tillTabOrderOnClickAddBookmarkButtonClick  TButtonRemoveSessionBookmarkButtonTagLeftTop)WidthSHeightAnchorsakTopakRight Caption&Ta bortTabOrderOnClickRemoveBookmarkButtonClick  TButtonUpSessionBookmarkButtonTag�LeftTop� WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickBookmarkButtonClick  TButtonDownSessionBookmarkButtonTagLeftTop� WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickBookmarkButtonClick   	TTabSheetSharedBookmarksSheetTagCaption   Delade bokmärken
ImageIndex
DesignSizez�   TListBoxSharedBookmarksListTagLeft
Top	WidthHeight� AnchorsakLeftakTopakRightakBottom DragModedmAutomatic
ItemHeightTabOrder OnClickBookmarksListClick
OnDblClickBookmarksListDblClick
OnDragDropBookmarksListDragDrop
OnDragOverBookmarksListDragOver	OnEndDragBookmarksListEndDrag	OnKeyDownBookmarksListKeyDownOnStartDragBookmarksListStartDrag  TButtonAddSharedBookmarkButtonTagLeftTop	WidthSHeightAnchorsakTopakRight Caption   &Lägg tillTabOrderOnClickAddBookmarkButtonClick  TButtonRemoveSharedBookmarkButtonTagLeftTop)WidthSHeightAnchorsakTopakRight Caption&Ta bortTabOrderOnClickRemoveBookmarkButtonClick  TButtonUpSharedBookmarkButtonTag�LeftTop� WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickBookmarkButtonClick  TButtonDownSharedBookmarkButtonTagLeftTop� WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickBookmarkButtonClick  TButtonShortCutSharedBookmarkButtonTagLeftTopIWidthSHeightAnchorsakTopakRight Caption   &Genväg...TabOrderOnClickShortCutBookmarkButtonClick    TButtonLocalDirectoryBrowseButtonLeft@TopWidthKHeightAnchorsakTopakRight Caption   Blädd&ra...TabOrderOnClickLocalDirectoryBrowseButtonClick  TButtonSwitchButtonLeftTop,WidthyHeightAnchorsakLeftakBottom CaptionP&latsprofiler...ModalResultTabOrderOnClickSwitchButtonClick  TButton
HelpButtonLeft@Top,WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick     TPF0TPreferencesDialogPreferencesDialogLeft�Top� HelpType	htKeywordHelpKeywordui_preferencesBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption   InställningarClientHeight�ClientWidth!Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize!� PixelsPerInch`
TextHeight TButtonOKButtonLeftTop�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCloseButtonLeftrTop�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TPanel	MainPanelLeft Top Width!Height�AlignalTopAnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneTabOrder  TPageControlPageControlLeft� Top Width�Height�
ActivePagePreferencesSheetAlignalClient	MultiLine	Style	tsButtonsTabOrderTabStopOnChangePageControlChange 	TTabSheetPreferencesSheetTagHelpType	htKeywordHelpKeywordui_pref_environmentCaption   Miljö
ImageIndex
TabVisible
DesignSize��  	TGroupBoxCommonPreferencesGroupLeftTopWidth�Height AnchorsakLeftakTopakRight Caption   BekräftelserTabOrder 
DesignSize�   	TCheckBoxConfirmOverwritingCheckLeftTop,WidtheHeightAnchorsakLeftakTopakRight Caption   &Överskrivning av filerTabOrderOnClickControlChange  	TCheckBoxConfirmDeletingCheckLeftTopCWidtheHeightAnchorsakLeftakTopakRight Caption%&Borttagning av filer (rekommenderad)TabOrderOnClickControlChange  	TCheckBoxConfirmClosingSessionCheckLeftTop� WidtheHeightAnchorsakLeftakTopakRight CaptionA&vsluta applikationenTabOrderOnClickControlChange  	TCheckBoxDDTransferConfirmationCheckLeftTop� WidtheHeightAnchorsakLeftakTopakRight Caption   D&ra && släpp-operationerTabOrderOnClickControlChange  	TCheckBoxContinueOnErrorCheckLeftTop� WidtheHeightAnchorsakLeftakTopakRight Caption*   Fortsätt vid &fel (avancerade användare)TabOrder	OnClickControlChange  	TCheckBoxConfirmExitOnCompletionCheckLeftTop� WidtheHeightAnchorsakLeftakTopakRight Caption.   Avsluta a&pplikationen vid slutförd operationTabOrderOnClickControlChange  	TCheckBoxConfirmResumeCheckLeftTopqWidtheHeightAnchorsakLeftakTopakRight Caption   &Återuppta överföringTabOrderOnClickControlChange  	TCheckBoxConfirmCommandSessionCheckLeftTop� WidtheHeightAnchorsakLeftakTopakRight Caption   Öppna separat &skalsessionTabOrderOnClickControlChange  	TCheckBoxConfirmRecyclingCheckLeftTopZWidtheHeightAnchorsakLeftakTopakRight Caption &Flytta filer till papperskorgenTabOrderOnClickControlChange  	TCheckBoxConfirmTransferringCheckLeftTopWidtheHeightAnchorsakLeftakTopakRight Caption   &Överföring av filerTabOrder OnClickControlChange   	TGroupBoxNotificationsGroupLeftTopWidth�HeightIAnchorsakLeftakTopakRight CaptionMeddelandenTabOrder
DesignSize�I  TLabelBeepOnFinishAfterTextLeftxTopWidthHeightAnchorsakTopakRight Captions  	TCheckBoxBeepOnFinishCheckLeftTopWidth$HeightAnchorsakLeftakTopakRight Caption=   S&ystemljud när operationen är klar, om den pågår mer änTabOrder OnClickControlChange  TUpDownEditBeepOnFinishAfterEditLeft:TopWidth9Height	AlignmenttaRightJustify	Increment       �@MaxValue      ��@AnchorsakTopakRight 	MaxLengthTabOrderOnChangeControlChange  	TCheckBoxBalloonNotificationsCheckLeftTop.WidthlHeightAnchorsakLeftakTopakRight CaptionK   Visa ballong&meddelanden i aktivitetsfältets statusområde (systemfältet)TabOrderOnClickControlChange    	TTabSheetLogSheetTagHelpType	htKeywordHelpKeywordui_pref_loggingCaptionLoggning
ImageIndex
TabVisible
DesignSize��  	TGroupBoxLoggingGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight Caption   Alternativ för loggningTabOrder 
DesignSize��   TLabelLogWindowLinesTextLeftGTop� WidthHeightAnchorsakTopakRight Captionrader  	TCheckBoxLogToFileCheckLeftTop/WidthgHeightAnchorsakLeftakTopakRight CaptionLogga till &fil:TabOrderOnClickControlChange  TFilenameEditLogFileNameEdit3Left(TopEWidthOHeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPathEditAfterDialog
DefaultExtlogFilter4Sessionsloggfilar (*.log)|*.log|Alla filer (*.*)|*.*DialogOptionsofHideReadOnlyofPathMustExist DialogTitle   Välj fil för sessionslogg.OnCreateEditDialogPathEditCreateEditDialogClickKey@AnchorsakLeftakTopakRight TabOrderTextLogFileNameEdit3OnChangeControlChange  	TCheckBoxLogShowWindowCheckLeftTopxWidthGHeightCaption   Visa loggf&önster:TabOrderOnClickControlChange  TRadioButtonLogWindowCompleteButtonLeft(Top� Width/HeightCaptionVisa &hela sessionenTabOrderOnClickControlChange  TRadioButtonLogWindowLinesButtonLeft(Top� Width� HeightAnchorsakLeftakTopakRight CaptionVisa endast &senasteTabOrderOnClickControlChange  TUpDownEditLogWindowLinesEditLeft� Top� WidthYHeight	AlignmenttaRightJustify	Increment       �@MaxValue      @�@MinValue       �@Value       �@AnchorsakTopakRight TabOrder	OnChangeControlChange  TPanelLogFilePanelLeft(Top]Width	HeightAnchorsakLeftakTopakRight 
BevelOuterbvNoneTabOrder TRadioButtonLogFileAppendButtonLeft TopWidthjHeightCaption   L&ägg tillTabOrder OnClickControlChange  TRadioButtonLogFileOverwriteButtonLeftpTopWidthjHeightCaption   Sk&riv överTabOrderOnClickControlChange   	TComboBoxLogProtocolComboLeft TopWidthwHeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChangeControlChangeItems.StringsNormalDebug 1Debug 2   TStaticTextLogFileNameHintTextLeft%Top[WidthRHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	   &mönsterTabOrderTabStop	  	TCheckBoxEnableLoggingCheckLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption!   Aktivera &sessionslogg på nivå:TabOrder OnClickControlChange   	TGroupBoxActionsLoggingGroupLeftTop� Width�HeightVAnchorsakLeftakTopakRight CaptionXML-loggTabOrder
DesignSize�V  TFilenameEditActionsLogFileNameEditLeft(Top+WidthOHeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPathEditAfterDialog
DefaultExtxmlFilter0XML-loggfiler (*.xml)|*.xml|Alla filer (*.*)|*.*DialogOptionsofHideReadOnlyofPathMustExist DialogTitle   Välj fil för XML-logg.OnCreateEditDialogPathEditCreateEditDialogClickKey@AnchorsakLeftakTopakRight TabOrderTextActionsLogFileNameEditOnChangeControlChange  TStaticTextActionsLogFileNameHintTextLeft%TopAWidthRHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	   möns&terTabOrderTabStop	  	TCheckBoxEnableActionsLoggingCheckLeftTopWidthgHeightAnchorsakLeftakTopakRight CaptionAktivera &XML-logg till fil:TabOrder OnClickControlChange    	TTabSheetGeneralSheetTagHelpType	htKeywordHelpKeywordui_pref_interfaceCaption   Gränssnitt
ImageIndex
TabVisible
DesignSize��  TLabelInterfaceChangeLabelLeftTopWidth� HeightCaption.   Ändringar kommer att gälla vid nästa start.  	TGroupBox
ThemeGroupLeftTop� Width�Height4AnchorsakLeftakTopakRight CaptionTemaTabOrder 
DesignSize�4  TLabelLabel7LeftTopWidthRHeightCaption   Gränssnitts&tema:FocusControl
ThemeCombo  	TComboBox
ThemeComboLeft� TopWidth� HeightStylecsDropDownListAnchorsakLeftakTopakRight TabOrder Items.StringsSystem	Office XPOffice 2003    	TGroupBoxInterfaceGroupLeftTopWidth�Height� AnchorsakLeftakTopakRightakBottom Caption   AnvändargränssnittTabOrder
DesignSize��   TLabelCommanderDescriptionLabel2Left� TopWidth� HeightsAnchorsakLeftakTopakRight AutoSizeCaption�   - två paneler (vänster för lokal katalog, höger för fjärrkatalog)
- snabbkommandon som i Norton Commander (och andra liknande program som Total Commander, Midnight Commander...)
- dra && släpp till/från båda panelernaWordWrap	OnClickCommanderClick  TLabelExplorerDescriptionLabelLeft� Top� Width� Height>AnchorsakLeftakTopakRight AutoSizeCaptionK   - endast fjärrkatalog
- snabbkommandon som i Utforskaren
- dra && släppWordWrap	OnClickExplorerClick  TImageCommanderInterfacePictureLeft7Top)Width Height AutoSize	Picture.Data
`  	TPngImage�PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?�@�Q��k^x�V���7?��׀9�VI#]m��S� t #�j6Qtu��#�P�v^Ɇ�<z���ڐ,'52|:я����Q:� Cw�Y�(Du���}$R6� CW�=Y�,Bu�{�>66@\W�@�!�@t&�3t��
�k�Y!+4�;t@�u�b�A��t$���;�8 �>h��Fw�ۣ�GA弃�I�D�t b��7Gz�B|^f��|�W�?�Кh���|�/`XF�Dm�Q�
�n�J��Z�� -�ɷ`q .}`�	�b�hxy���`�]p��j �@�/�2|� �	�qAY��CS���H�q�4@e�G���]	���a�t�,�gP
���jPc�-D~�a0�k�"㪩�����A�J٣9�������F�E�PI��xz���o�5�dQ�^�a�i�a��X[�~��B$}�������0�y	������˃�}�P�#8-���Ӳ���x����`lZT5+�|rNhx�����%�#��J�r@��#��6�Ba�u=^���Q@w�����.C��q@�2�AYe��'B�u@�2�QP	ի���{�G��s����D�:Pr)Cu��=]$�	t@9)@�+�Ғ���	�`�܍��	)Ti�R�W�b��S����@�w  G��Ш���    IEND�B`�OnClickCommanderClick  TImageExplorerInterfacePictureLeft7Top� Width Height AutoSize	Picture.Data
L  	TPngImage�PNG

   IHDR           szz�   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?�@F�x̋�12�W�����=կ�Sh7�����J��i=�_NM`$�j6QTw��#ˈw��yTw@pR�r���}Tw��u�xu�,�c�4���,?�U���Zm(rs�N��S����m1�x~�,�������E÷K�p6�^3�ܤӭpv�i5���+!�O@�P�p@C+��/���l�&��C��)�����	x�����@Ω�x��q@��#p�Q6v���_����@�䗓}Jp��݅U��k�J��'������B5�rZ��(����?�%��1hz�3Ъ�Bq��m`�;��e�K1�xU����B0i�-��� 5=�
Z��(8���BC�JX)�����ɻ>�ٹn(r�JWP)��3!���\q����%���V��@��'pv�����TJ�8��Բ��`�$���Wހ�+�5P��t��pj�Ѫ��;��gi��cV���D	��Ip �R� *a�v �R� *a�v ��d^:.�7:E�]D[�2j[�tP	K�`�$Ӵ����uL7�rꨕz�
��h�JI�vD��_%j���U�����(r�+�JX������JX����D�ʁJX������JX��mVH��+�I6�  ����,Md    IEND�B`�Transparent	OnClickExplorerClick  TRadioButtonCommanderInterfaceButton2LeftTopWidthtHeightCaption
&CommanderChecked	TabOrder TabStop	OnClickControlChange  TRadioButtonExplorerInterfaceButton2LeftTop� WidthoHeightCaption&UtforskareTabOrderOnClickControlChange    	TTabSheetPanelsSheetTagHelpType	htKeywordHelpKeywordui_pref_panelsCaptionPaneler
ImageIndex
TabVisible
DesignSize��  	TGroupBoxPanelsCommonGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight Caption   AllmäntTabOrder 
DesignSize��   	TCheckBoxShowHiddenFilesCheckLeftTopWidtheHeightAnchorsakLeftakTopakRight CaptionVi&sa dolda filer (CTRL+ALT+H)TabOrder OnClickControlChange  	TCheckBoxDefaultDirIsHomeCheckLeftTopEWidtheHeightAnchorsakLeftakTopakRight Caption!   Standardkatalog är &hemkatalogenTabOrderOnClickControlChange  	TCheckBoxDeleteToRecycleBinCheckLeftTop-WidtheHeightAnchorsakLeftakTopakRight Caption'Ta bort lokala filer till papperskorgenTabOrderOnClickControlChange  	TCheckBoxPreservePanelStateCheckLeftTop]WidtheHeightAnchorsakLeftakTopakRight Caption4   Kom i&håg panelens' tillstånd när session växlasTabOrderOnClickControlChange  	TCheckBoxRenameWholeNameCheckLeftTopuWidtheHeightAnchorsakLeftakTopakRight Caption&   Välj &hela namnet när filen döps omTabOrderOnClickControlChange  	TCheckBoxFormatSizeBytesCheckLeftTop� WidtheHeightAnchorsakLeftakTopakRight Caption Visa filstorlekar i kort &formatTabOrderOnClickControlChange  	TCheckBoxFullRowSelectCheckLeftTop� WidtheHeightAnchorsakLeftakTopakRight Caption   Välja med h&ela radenTabOrderOnClickControlChange   	TGroupBoxDoubleClickGroupLeftTop� Width�HeightJAnchorsakLeftakTopakRight CaptionDubbelklickTabOrder
DesignSize�J  TLabelDoubleClickActionLabelLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption'   &Operation att utföra vid dubbelklick:FocusControlDoubleClickActionCombo  	TCheckBox"CopyOnDoubleClickConfirmationCheckLeft Top-WidthTHeightAnchorsakLeftakTopakRight Caption+   &Bekräfta kopiera vid dubbelklickoperationTabOrderOnClickControlChange  	TComboBoxDoubleClickActionComboLeftTopWidthlHeightStylecsDropDownListAnchorsakTopakRight TabOrder OnChangeControlChangeItems.Strings   ÖppnaKopieraRedigera     	TTabSheetCommanderSheetTagHelpType	htKeywordHelpKeywordui_pref_commanderCaption	Commander
ImageIndex
TabVisible
DesignSize��  TLabelLabel3LeftTopWidth�HeightAnchorsakLeftakTopakRight AutoSizeCaptionV   Inställningar på den här fliken gäller endast för Norton Commander-gränssnittet.WordWrap	  	TGroupBoxPanelsGroupLeftTop&Width�HeightcAnchorsakLeftakTopakRight CaptionPanelerTabOrder 
DesignSize�c  TLabelLabel8LeftTopWidthtHeightCaptionVal av &utforskarstil:FocusControlNortonLikeModeCombo  	TCheckBoxSwappedPanelsCheckLeftTop-WidtheHeightAnchorsakLeftakTopakRight Caption6   B&yt paneler (lokal till höger, fjärr till vänster)TabOrderOnClickControlChange  	TComboBoxNortonLikeModeComboLeft� TopWidth� HeightStylecsDropDownListAnchorsakLeftakTopakRight TabOrder OnChangeControlChangeItems.StringsAldrigBara musMus och tangentbord   	TCheckBoxTreeOnLeftCheckLeftTopEWidtheHeightAnchorsakLeftakTopakRight Caption(   Visa &katalogträd vänster om fillistanTabOrderOnClickControlChange   	TGroupBoxCommanderMiscGroupLeftTop� Width�HeightMAnchorsakLeftakTopakRight Caption   ÖvrigtTabOrder
DesignSize�M  TLabelLabel10LeftTopWidth^HeightCaption&KortkommandonFocusControlExplorerKeyboardShortcutsCombo  	TCheckBoxUseLocationProfilesCheckLeftTop-WidtheHeightAnchorsakLeftakTopakRight Caption7   &Använd platsprofiler istället för katalogbokmärkenTabOrderOnClickControlChange  	TComboBoxExplorerKeyboardShortcutsComboLeft� TopWidth� HeightStylecsDropDownListAnchorsakLeftakTopakRight TabOrder OnChangeControlChangeItems.Strings	CommanderUtforskaren    	TGroupBoxCompareCriterionsGroupLeftTop� Width�HeightJAnchorsakLeftakTopakRight Caption   Jämför katalogkriteriumTabOrder
DesignSize�J  	TCheckBoxCompareByTimeCheckLeftTopWidtheHeightAnchorsakLeftakTopakRight Caption   Jämför efter &tidTabOrder OnClickControlChange  	TCheckBoxCompareBySizeCheckLeftTop-WidtheHeightAnchorsakLeftakTopakRight Caption   Jämför efter &storlekTabOrderOnClickControlChange    	TTabSheetExplorerSheetTagHelpType	htKeywordHelpKeywordui_pref_explorerCaptionUtforskaren
ImageIndex
TabVisible
DesignSize��  TLabelLabel4LeftTopWidth�HeightAnchorsakLeftakTopakRight AutoSizeCaptionM   Inställningar på den här fliken gäller endast för utforskargränssnittetWordWrap	  	TGroupBox	GroupBox2LeftTop&Width�Height6AnchorsakLeftakTopakRight CaptionVisaTabOrder 
DesignSize�6  	TCheckBoxShowFullAddressCheckLeftTopWidtheHeightAnchorsakLeftakTopakRight Caption2   Vi&sa den fullständiga sökvägen i adressfältetTabOrder OnClickControlChange    	TTabSheetEditorSheetTagHelpType	htKeywordHelpKeywordui_pref_editorCaptionEditor
ImageIndex
TabVisible
DesignSize��  	TGroupBoxInternalEditorGroupLeftTop� Width�Height� AnchorsakLeftakRightakBottom Caption   Alternativ för intern editorTabOrder
DesignSize��   TLabelEditorFontLabelLeft� Top1Width� HeightXAnchorsakTopakRight AutoSizeCaptionEditorFontLabelColor	clBtnFaceParentColorTransparent
OnDblClickEditorFontLabelDblClick  TLabelLabel9LeftTop/WidthGHeightCaption&Tabulatorstorlek:FocusControlEditorTabSizeEdit  TLabelLabel11LeftTop_WidthUHeightCaptionStandard&kodning:FocusControlEditorEncodingCombo  TButtonEditorFontButtonLeft� TopWidthiHeightAnchorsakTopakRight Caption   &Välj font...TabOrderOnClickEditorFontButtonClick  	TCheckBoxEditorWordWrapCheckLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption   Ko&rta av långa raderTabOrder OnClickControlChange  TUpDownEditEditorTabSizeEditLeftTop@Width� Height	AlignmenttaRightJustifyMaxValue       �@MinValue       ��?Value       ��?AnchorsakLeftakTopakRight 	MaxLengthTabOrderOnChangeControlChange  	TComboBoxEditorEncodingComboLeftToppWidth� HeightStylecsDropDownListAnchorsakLeftakTopakRight 	MaxLengthTabOrderOnChangeControlChange   	TGroupBoxEditorPreferenceGroupLeftTopWidth�Height� AnchorsakLeftakTopakRightakBottom Caption   EditorinställningarTabOrder 
DesignSize��   	TListViewEditorListView3LeftTopWidthdHeight� AnchorsakLeftakTopakRightakBottom ColumnsCaptionEditorWidth�  CaptionMaskWidthF CaptionTextTagWidth-  ColumnClickDoubleBuffered	DragModedmAutomaticHideSelection	OwnerData	ReadOnly		RowSelect	ParentDoubleBufferedTabOrder 	ViewStylevsReportOnDataEditorListView3Data
OnDblClickEditorListView3DblClick	OnEndDragListViewEndDrag
OnDragDropEditorListView3DragDrop
OnDragOverListViewDragOver	OnKeyDownEditorListView3KeyDownOnSelectItemListViewSelectItemOnStartDragListViewStartDrag  TButtonAddEditorButtonLeftTop� WidthSHeightAnchorsakLeftakBottom Caption   &Lägg till...TabOrderOnClickAddEditEditorButtonClick  TButtonEditEditorButtonLeftpTop� WidthSHeightAnchorsakLeftakBottom Caption&Redigera...TabOrderOnClickAddEditEditorButtonClick  TButtonUpEditorButtonLeft"Top� WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickUpDownEditorButtonClick  TButtonDownEditorButtonLeft"Top� WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickUpDownEditorButtonClick  TButtonRemoveEditorButtonLeftTop� WidthSHeightAnchorsakLeftakBottom Caption&Ta bortTabOrderOnClickRemoveEditorButtonClick    	TTabSheetIntegrationSheetTag	HelpType	htKeywordHelpKeywordui_pref_integrationCaptionIntegrering
ImageIndex
TabVisible
DesignSize��  	TGroupBoxShellIconsGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight CaptionWindowsskalTabOrder 
DesignSize��   TButtonDesktopIconButtonLeftTopWidtheHeightAnchorsakLeftakTopakRight Caption   Skapa en ikon på skrivbor&detTabOrder OnClickIconButtonClick  TButtonQuickLaunchIconButtonLeftTop8WidtheHeightAnchorsakLeftakTopakRight CaptionSkapa en sna&bbstartsikonTabOrderOnClickIconButtonClick  TButtonSendToHookButtonLeftTopXWidtheHeightAnchorsakLeftakTopakRight CaptionB   Skapa genväg för överföring i utforskarens '&Skicka till'-menyTabOrderOnClickIconButtonClick  TButtonRegisterAsUrlHandlersButtonLeftTop� WidtheHeightAnchorsakLeftakTopakRight Caption)   Registrera för att hantera &URL-adresserTabOrderOnClick RegisterAsUrlHandlersButtonClick  TButtonAddSearchPathButtonLeftTop� WidtheHeightAnchorsakLeftakTopakRight Caption7   Lägg till sökvägen till WinSCP i miljövaribeln PATHTabOrderOnClickAddSearchPathButtonClick  TStaticTextShellIconsText2Left+ToptWidthJHeightHint   För att lägga till genvägar, som direkt öppnar webbplats, använd ikonkommandon i 'Hantera'-menyn i dialogrutan inloggning.	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaptionAssociera ikoner med webbplatsTabOrderTabStop	    	TTabSheetCustomCommandsSheetTag
HelpType	htKeywordHelpKeywordui_pref_commandsCaption	Kommandon
ImageIndex	
TabVisible
DesignSize��  	TGroupBoxCustomCommandsGroupLeftTopWidth�HeightvAnchorsakLeftakTopakRightakBottom CaptionEgna kommandonTabOrder 
DesignSize�v  	TListViewCustomCommandsViewLeftTopWidthdHeight
AnchorsakLeftakTopakRightakBottom ColumnsCaptionBeskrivningWidthU CaptionKommandoWidth�  CaptionL/FTagWidth# CaptionK/RTagWidth(  ColumnClickDoubleBuffered	DragModedmAutomaticHideSelection	OwnerData	ReadOnly		RowSelect	ParentDoubleBufferedTabOrder 	ViewStylevsReportOnDataCustomCommandsViewData
OnDblClickCustomCommandsViewDblClick	OnEndDragListViewEndDrag
OnDragDropCustomCommandsViewDragDrop
OnDragOverListViewDragOver	OnKeyDownCustomCommandsViewKeyDownOnSelectItemListViewSelectItemOnStartDragListViewStartDrag  TButtonAddCommandButtonLeftTop-WidthSHeightAnchorsakLeftakBottom Caption   &Lägg till...TabOrderOnClickAddEditCommandButtonClick  TButtonRemoveCommandButtonLeftTopMWidthSHeightAnchorsakLeftakBottom Caption&Ta bortTabOrderOnClickRemoveCommandButtonClick  TButtonUpCommandButtonLeft"Top-WidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickUpDownCommandButtonClick  TButtonDownCommandButtonLeft"TopMWidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickUpDownCommandButtonClick  TButtonEditCommandButtonLeftpTop-WidthSHeightAnchorsakLeftakBottom Caption&Redigera...TabOrderOnClickAddEditCommandButtonClick    	TTabSheetDragDropSheetTagHelpType	htKeywordHelpKeywordui_pref_dragdropCaption   Dra & släpp
ImageIndex

TabVisible
DesignSize��  	TGroupBoxDragDropDownloadsGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight Caption   Dra && släpp nerladdningarTabOrder 
DesignSize��   TLabelDDExtEnabledLabelLeft#TopDWidthYHeight5AnchorsakLeftakTopakRight AutoSizeCaption�   Möjliggör direkt nerladdningar till vanliga lokala kataloger (t. ex. utforskaren). Tillåter inte nerladdningar till andra destinationer (ZIP-arkiv, FTP, etc.)WordWrap	OnClickDDExtLabelClick  TLabelDDExtDisabledLabelLeft#Top� WidthZHeight6AnchorsakLeftakTopakRight AutoSizeCaption�   Möjliggör nerladdningar till valfri destination (vanliga kataloger, ZIP-arkiv, FTP, etc.). Filer laddas först ner till en temporär katalog och flyttas därefter till destinationen.WordWrap	OnClickDDExtLabelClick  TRadioButtonDDExtEnabledButtonLeftTop0WidthlHeightAnchorsakLeftakTopakRight Caption   Använd &skaltilläggTabOrderOnClickControlChange  TRadioButtonDDExtDisabledButtonLeftTop|WidthdHeightAnchorsakLeftakTopakRight Caption   Använd &temporär katalogTabOrderOnClickControlChange  TPanelDDExtDisabledPanelLeft"Top� Width;Height3
BevelOuterbvNoneTabOrder
DesignSize;3  	TCheckBoxDDWarnLackOfTempSpaceCheckLeft TopWidth;HeightAnchorsakLeftakTopakRight Caption)   &Varna vid otillräckligt med diskutrymmeTabOrder OnClickControlChange  	TCheckBoxDDWarnOnMoveCheckLeft TopWidth;HeightAnchorsakLeftakTopakRight Caption&   Varna vid &flytt via temporär katalogTabOrderOnClickControlChange   	TCheckBoxDDAllowMoveInitCheckLeftTopWidthlHeightAnchorsakLeftakTopakRight Caption?   Tillåt f&lyttning från fjärrkatalog till andra applikationerTabOrder OnClickControlChange    	TTabSheet
QueueSheetTagHelpType	htKeywordHelpKeywordui_pref_backgroundCaptionBakgrund
ImageIndex
TabVisible
DesignSize��  	TGroupBox
QueueGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight Caption   Överföringar i bakgrundenTabOrder 
DesignSize��   TLabelLabel5LeftTopWidth� HeightCaption)   &Maximalt antal samtidiga överföringar:FocusControlQueueTransferLimitEdit  TLabelQueueKeepDoneItemsCheckLeftTop� Width� HeightCaption*   Visa avslutade överföringar i kön för:FocusControlQueueKeepDoneItemsForComboOnClickControlChange  TUpDownEditQueueTransferLimitEditLeft0TopWidthIHeight	AlignmenttaRightJustifyMaxValue       �@MinValue       ��?Value       ��?AnchorsakTopakRight 	MaxLengthTabOrder   	TCheckBoxQueueAutoPopupCheckLeftTop� WidthqHeightAnchorsakLeftakTopakRight CaptionC   Visa bakgrundsöverföringarnas prompt &automatiskt vid inaktivitetTabOrder  	TCheckBox
QueueCheckLeftTopJWidthqHeightAnchorsakLeftakTopakRight Caption$   &Överför som standard i bakgrundenTabOrder  	TCheckBoxQueueNoConfirmationCheckLeftTopzWidthqHeightAnchorsakLeftakTopakRight Caption1   I&ngen bekräftelser för bakgrundsöverföringarTabOrder  	TCheckBoxQueueIndividuallyCheckLeftTopbWidthqHeightAnchorsakLeftakTopakRight Caption/   &Lägg till varje fil individuellt som standardTabOrder  	TCheckBoxEnableQueueByDefaultCheckLeftTop2WidthqHeightAnchorsakLeftakTopakRight Caption$   &Aktivera köbehandling som standardTabOrder  	TComboBoxQueueKeepDoneItemsForComboLeftTop� WidthaHeightStylecsDropDownListAnchorsakTopakRight 	MaxLengthTabOrderOnChangeControlChangeItems.StringsAldrig15 sekunder1 minut
15 minuter1 timmeAlltid    	TGroupBoxQueueViewGroupLeftTop� Width�HeightcAnchorsakLeftakTopakRight Caption   KölistaTabOrder
DesignSize�c  TRadioButtonQueueViewShowButtonLeftTopWidthqHeightAnchorsakLeftakTopakRight CaptionVi&saTabOrder   TRadioButtonQueueViewHideWhenEmptyButtonLeftTop-WidthqHeightAnchorsakLeftakTopakRight Caption   &Dölj ifall tomTabOrder  TRadioButtonQueueViewHideButtonLeftTopEWidthqHeightAnchorsakLeftakTopakRight Caption   &DöljTabOrder    	TTabSheetStorageSheetTagHelpType	htKeywordHelpKeywordui_pref_storageCaptionLagring
ImageIndex
TabVisible
DesignSize��  	TGroupBoxStorageGroupLeftTopWidth�HeightHAnchorsakLeftakTopakRight Caption   Inställningar för lagringTabOrder 
DesignSize�H  TRadioButtonRegistryStorageButtonLeftTopWidthhHeightAnchorsakLeftakTopakRight CaptionWindowsre&gistretTabOrder OnClickControlChange  TRadioButtonIniFileStorageButton2LeftTop-WidthhHeightAnchorsakLeftakTopakRight Caption&INI-fil (winscp.ini)TabOrderOnClickControlChange   	TGroupBoxTemporaryDirectoryGrouoLeftTopXWidth�Height� AnchorsakLeftakTopakRight Caption   Temporär katalogTabOrder
DesignSize��   TLabelLabel6LeftTopWidthhHeightAnchorsakLeftakTopakRight AutoSizeCaption?   Ange var nerladdade och redigerade filer ska sparas temporärt.WordWrap	  TRadioButton DDSystemTemporaryDirectoryButtonLeftTop-WidthhHeightAnchorsakLeftakTopakRight Caption%   &Använd systemets temporära katalogTabOrder OnClickControlChange  TRadioButton DDCustomTemporaryDirectoryButtonLeftTopEWidth� HeightCaption   Använd den här &katalogen:TabOrderOnClickControlChange  TDirectoryEditDDTemporaryDirectoryEditLeft� TopAWidth� HeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPathEditAfterDialog
DialogText2   Välj katalog för temporära dra && släpp filer.ClickKey@AnchorsakLeftakTopakRight TabOrderTextDDTemporaryDirectoryEditOnClickControlChange  	TCheckBoxTemporaryDirectoryCleanupCheckLeftTop� WidthhHeightAnchorsakLeftakTopakRight Caption.   &Rensa gamla temporära kataloger vid uppstartTabOrderOnClickControlChange  	TCheckBox%ConfirmTemporaryDirectoryCleanupCheckLeft Top� WidthXHeightAnchorsakLeftakTopakRight Caption   &Fråga innan rensningTabOrderOnClickControlChange  	TCheckBox$TemporaryDirectoryAppendSessionCheckLeftTop^WidthhHeightAnchorsakLeftakTopakRight Caption3   Lägg till &sessionsnamn till temporära sökvägenTabOrderOnClickControlChange  	TCheckBox!TemporaryDirectoryAppendPathCheckLeftTopwWidthhHeightAnchorsakLeftakTopakRight Caption5   Lägg till f&järrsökväg till temporära sökvägenTabOrderOnClickControlChange   	TGroupBoxOtherStorageGroupLeftTop%Width�Height5AnchorsakLeftakTopakRight Caption   ÖvrigtTabOrder
DesignSize�5  TLabelRandomSeedFileLabelLeftTopWidthVHeightCaption   Sl&umptalsfröfil:FocusControlRandomSeedFileEdit  TFilenameEditRandomSeedFileEditLeft� TopWidth� HeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPathEditAfterDialog
DefaultExtlogFilter4   Slumptalsfröfiler (*.rnd|*.rnd|Alla filer (*.*)|*.*DialogOptionsofHideReadOnlyofPathMustExist DialogTitle   Välj fil för slumptalsfröOnCreateEditDialogPathEditCreateEditDialogClickKey@AnchorsakLeftakTopakRight TabOrder TextRandomSeedFileEditOnChangeControlChange    	TTabSheetTransferEnduranceSheetTagHelpType	htKeywordHelpKeywordui_pref_resumeCaptionTolerans
ImageIndex
TabVisible
DesignSize��  	TGroupBox	ResumeBoxLeftTopWidth�Height{AnchorsakLeftakTopakRight Caption@   Aktivera överföringspaus/överför till temporär filnamn förTabOrder  TLabelResumeThresholdUnitLabelLeft� TopGWidthHeightCaptionkBFocusControlResumeThresholdEdit  TRadioButtonResumeOnButtonLeftTopWidthIHeightCaptionA&lla filerTabOrder OnClickControlChange  TRadioButtonResumeSmartButtonLeftTop-Width� HeightCaption   Filer stö&rre än:TabOrderOnClickControlChange  TRadioButtonResumeOffButtonLeftTop]WidthIHeightCaptionA&vaktiveraTabOrderOnClickControlChange  TUpDownEditResumeThresholdEditLeft-TopCWidthTHeight	AlignmenttaRightJustify	Increment       �@MaxValue       �@TabOrderOnClickControlChange   	TGroupBoxSessionReopenGroupLeftTop� Width�Height� AnchorsakLeftakTopakRight Caption   Automatisk återanslutningTabOrder TLabelSessionReopenAutoLabelLeft"Top0WidthRHeightCaption   &Återanslut efter:FocusControlSessionReopenAutoEdit  TLabelSessionReopenAutoSecLabelLeftTop0Width'HeightCaptionsekunderFocusControlSessionReopenAutoEdit  TLabelSessionReopenTimeoutLabelLeftTop� WidthnHeightCaption   &Fortsätt återansluta i:FocusControlSessionReopenTimeoutEdit  TLabelSessionReopenTimeoutSecLabelLeftTop� Width'HeightCaptionsekunderFocusControlSessionReopenTimeoutEdit  TLabelSessionReopenAutoStallLabelLeft"Top� WidthRHeightCaption   Å&teranslut efter:FocusControlSessionReopenAutoStallEdit  TLabelSessionReopenAutoStallSecLabelLeftTop� Width'HeightCaptionsekunderFocusControlSessionReopenAutoStallEdit  TLabelSessionReopenAutoIdleLabelLeft"TopcWidthRHeightCaption   Å&teranslut efter:FocusControlSessionReopenAutoIdleEdit  TLabelSessionReopenAutoIdleSecLabelLeftTopcWidth'HeightCaptionsekunderFocusControlSessionReopenAutoIdleEdit  	TCheckBoxSessionReopenAutoCheckLeftTopWidthQHeightCaptionA   &Automatiskt återanslut session, om den bryts under överföringTabOrder OnClickControlChange  TUpDownEditSessionReopenAutoEditLeft� Top+WidthaHeight	AlignmenttaRightJustify	Increment       �@MaxValue       �@MinValue       ��?Value       �@	MaxLengthTabOrder  	TCheckBoxSessionReopenAutoIdleCheckLeftTopHWidthQHeightCaption9   Automatiskt återanslut session, om den &bryts under idleTabOrderOnClickControlChange  TUpDownEditSessionReopenTimeoutEditLeft� Top� WidthaHeight	AlignmenttaRightJustify	Increment       �@MaxValue      ��@	MaxLengthTabOrder
OnGetValue SessionReopenTimeoutEditGetValue
OnSetValue SessionReopenTimeoutEditSetValue  	TCheckBoxSessionReopenAutoStallCheckLeftTopzWidthQHeightCaption0   Automatiskt återanslut session, om den &stannarTabOrderOnClickControlChange  TUpDownEditSessionReopenAutoStallEditLeft� Top� WidthaHeight	AlignmenttaRightJustify	Increment       �@MaxValue       �@MinValue       ��?Value       �@	MaxLengthTabOrder  TUpDownEditSessionReopenAutoIdleEditLeft� Top^WidthaHeight	AlignmenttaRightJustify	Increment       �@MaxValue       �@MinValue       ��?Value       �@	MaxLengthTabOrder    	TTabSheetUpdatesSheetTagHelpType	htKeywordHelpKeywordui_pref_updatesCaptionUppdateringar
ImageIndex
TabVisible
DesignSize��  	TGroupBoxUpdatesGroupLeftTopWidth�Height3AnchorsakLeftakTopakRight Caption1Kontrollera automatisk om det finns uppdateringarTabOrder 
DesignSize�3  TLabelLabel12LeftTopWidthsHeightCaptionAutomatisk kontroll&period:FocusControlUpdatesPeriodCombo  	TComboBoxUpdatesPeriodComboLeftTopWidthbHeightStylecsDropDownListAnchorsakTopakRight TabOrder Items.StringsAldrigDagligVeckovis
   Månadsvis    	TGroupBoxUpdatesProxyGroupLeftTop� Width�Height� AnchorsakLeftakTopakRight Caption
AnslutningTabOrder
DesignSize��   TLabelUpdatesProxyHostLabelLeft"Top[WidthUHeightCaption   Proxy &värdnamn:FocusControlUpdatesProxyHostEdit  TLabelUpdatesProxyPortLabelLeftTop[Width?HeightAnchorsakTopakRight CaptionPo&rtnummer:FocusControlUpdatesProxyPortEdit  TUpDownEditUpdatesProxyPortEditLeftToplWidthbHeight	AlignmenttaRightJustifyMaxValue      ��@MinValue       ��?Value       ��?AnchorsakTopakRight TabOrder  TEditUpdatesProxyHostEditLeft"ToplWidth� HeightAnchorsakLeftakTopakRight 	MaxLength2TabOrderTextUpdatesProxyHostEdit  TRadioButtonUpdatesProxyCheckLeftTopEWidthmHeightAnchorsakLeftakTopakRight Caption   A&nvänd proxyserverTabOrderOnClickControlChange  TRadioButtonUpdatesDirectCheckLeftTopWidthmHeightAnchorsakLeftakTopakRight CaptionIngen &proxyTabOrder OnClickControlChange  TRadioButtonUpdatesAutoCheckLeftTop-WidthmHeightAnchorsakLeftakTopakRight Caption)   Detektera &automatisk proxyinställningarTabOrderOnClickControlChange   	TGroupBoxUpdatesOptionsGroupLeftTopAWidth�HeightQAnchorsakLeftakTopakRight Caption
AlternativTabOrder
DesignSize�Q  TLabelUpdatesBetaVersionsLabelLeftTopWidthvHeightCaption+Kontrollera ifall det finns &betaversioner:FocusControlUpdatesBetaVersionsCombo  	TComboBoxUpdatesBetaVersionsComboLeftTopWidthbHeightStylecsDropDownListAnchorsakTopakRight TabOrder   	TCheckBoxCollectUsageCheckLeftTop1WidthHeightAnchorsakLeftakTopakRight Caption"   Tillåt &anonym användarstatistikTabOrderOnClickControlChange  TButtonUsageViewButtonLeftTop-WidthbHeightAnchorsakTopakRight CaptionVisa &statistikTabOrderOnClickUsageViewButtonClick    	TTabSheetCopyParamListSheetTagHelpType	htKeywordHelpKeywordui_pref_presetsCaption	   Överför
ImageIndex
TabVisible
DesignSize��  	TGroupBoxCopyParamListGroupLeftTopWidth�HeightvAnchorsakLeftakTopakRightakBottom Caption   Överför förinställningarTabOrder 
DesignSize�v  TLabelCopyParamLabelLeftTop� WidthbHeight5AnchorsakLeftakRightakBottom AutoSizeCaptionCopyParamLabelWordWrap	OnClickCopyParamLabelClick  	TListViewCopyParamListViewLeftTopWidthdHeight� AnchorsakLeftakTopakRightakBottom ColumnsCaption   Beskrivning förinställningarWidthd Caption
AutomatiskTagWidth(  ColumnClickDoubleBuffered	DragModedmAutomaticHideSelection	OwnerData	ReadOnly		RowSelect	ParentDoubleBufferedTabOrder 	ViewStylevsReportOnCustomDrawItemCopyParamListViewCustomDrawItemOnDataCopyParamListViewData
OnDblClickCopyParamListViewDblClick	OnEndDragListViewEndDrag
OnDragDropCopyParamListViewDragDrop
OnDragOverListViewDragOver	OnKeyDownCopyParamListViewKeyDownOnSelectItemListViewSelectItemOnStartDragListViewStartDrag  TButtonAddCopyParamButtonLeftTopWidthSHeightAnchorsakLeftakBottom Caption   &Lägg till...TabOrderOnClickAddCopyParamButtonClick  TButtonRemoveCopyParamButtonLeftTop9WidthSHeightAnchorsakLeftakBottom Caption&Ta bortTabOrderOnClickRemoveCopyParamButtonClick  TButtonUpCopyParamButtonLeft!TopWidthSHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickUpDownCopyParamButtonClick  TButtonDownCopyParamButtonLeft!Top9WidthSHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickUpDownCopyParamButtonClick  TButtonEditCopyParamButtonLeftpTopWidthSHeightAnchorsakLeftakBottom Caption&Redigera...TabOrderOnClickEditCopyParamButtonClick  TButtonDuplicateCopyParamButtonLeftpTop9WidthSHeightAnchorsakLeftakBottom Caption&Dubblera...TabOrderOnClickDuplicateCopyParamButtonClick  	TCheckBoxCopyParamAutoSelectNoticeCheckLeftTopXWidthbHeightAnchorsakLeftakRightakBottom CaptionS   &Meddela när överföringsinställningarna automatiskt använder de förinställdaTabOrderOnClickControlChange    	TTabSheetWindowSheetTagHelpType	htKeywordHelpKeywordui_pref_windowCaption   Fönster
ImageIndex
TabVisible
DesignSize��  	TGroupBoxPathInCaptionGroupLeftTop� Width�Height^AnchorsakLeftakTopakRight Caption   Sökväg i fönstertitelTabOrder
DesignSize�^  TRadioButtonPathInCaptionFullButtonLeftTopWidthiHeightAnchorsakLeftakTopakRight Caption   Visa &lång sökvägTabOrder   TRadioButtonPathInCaptionShortButtonLeftTop,WidthiHeightAnchorsakLeftakTopakRight Caption   Visa &kort sökvägTabOrder  TRadioButtonPathInCaptionNoneButtonLeftTopCWidthiHeightAnchorsakLeftakTopakRight Caption
Visa &inteTabOrder   	TGroupBoxWindowMiscellaneousGroupLeftTop� Width�Height5AnchorsakLeftakTopakRight Caption   ÖvrigtTabOrder
DesignSize�5  	TCheckBoxMinimizeToTrayCheckLeftTopWidthiHeightAnchorsakLeftakTopakRight CaptionN   &Minimera huvudfönstret till aktivitetsfältets statusområde (systemfältet)TabOrder OnClickControlChange   	TGroupBoxWorkspacesGroupLeftTopWidth�HeightuAnchorsakLeftakTopakRight Caption
ArbetsytorTabOrder 
DesignSize�u  TLabelAutoWorkspaceLabelLeft-Top-WidthzHeightCaption&Standardnamn arbetsyta:FocusControlAutoWorkspaceCombo  	TCheckBoxAutoSaveWorkspaceCheckLeftTopWidthiHeightAnchorsakLeftakTopakRight Caption'Spara &automatiskt arbetsyta vid avslutTabOrder OnClickControlChange  	TComboBoxAutoWorkspaceComboLeft-Top=WidthLHeightAnchorsakLeftakTopakRight DropDownCountTabOrderOnClickControlChange  	TCheckBoxAutoSaveWorkspacePasswordsCheckLeft-TopWWidthLHeightAnchorsakLeftakTopakRight Caption#Save &passwords (not recommended) XTabOrderOnClickControlChange    	TTabSheetSecuritySheetTagHelpType	htKeywordHelpKeywordui_pref_securityCaption	   Säkerhet
ImageIndex
TabVisible
DesignSize��  	TGroupBoxMasterPasswordGroupLeftTopWidth�Height\AnchorsakLeftakTopakRight Caption   HuvudlösenordTabOrder 
DesignSize�\  TButtonSetMasterPasswordButtonLeftTop3WidtheHeightAnchorsakLeftakTopakRight Caption   Ä&ndra huvudlösenord...TabOrderOnClickSetMasterPasswordButtonClick  	TCheckBoxUseMasterPasswordCheckLeftTopWidthdHeightAnchorsakLeftakTopakRight Caption   An&vänd huvudlösenordTabOrder OnClickUseMasterPasswordCheckClick   	TGroupBoxPasswordGroupBoxLeftTopjWidth�Height4AnchorsakLeftakTopakRight Caption   SessionslösenordTabOrder
DesignSize�4  	TCheckBoxSessionRememberPasswordCheckLeftTopWidthdHeightAnchorsakLeftakTopakRight Caption1   Kom ihåg &lösenord under sessionens varaktighetTabOrder     	TTabSheetIntegrationAppSheetTagHelpType	htKeywordHelpKeywordui_pref_integration_appCaptionApplikationer
ImageIndex
TabVisible
DesignSize��  	TGroupBoxExternalAppsGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight CaptionExterna applikationerTabOrder 
DesignSize��   TLabelPuttyPathLabelLeftTopWidth� HeightCaption    &PuTTY/Terminal klient sökväg:FocusControlPuttyPathEdit  TLabelPuttyRegistryStorageKeyLabelLeftTop� Width^HeightCaptionPuTTY registernyc&kelFocusControlPuttyRegistryStorageKeyEdit  THistoryComboBoxPuttyPathEditLeftTop&WidthHeightAnchorsakLeftakTopakRight TabOrder OnChangePuttyPathEditChange  	TCheckBoxPuttyPasswordCheck2LeftTopSWidthaHeightAnchorsakLeftakTopakRight Caption?   &Kom ihåg sessionslösenord och överför det till PuTTY (SSH)TabOrder  	TCheckBoxAutoOpenInPuttyCheckLeftTop� WidthaHeightAnchorsakLeftakTopakRight Caption)   &Öppna automatiskt en ny session i PuTTYTabOrder  TButtonPuttyPathBrowseButtonLeft/Top$WidthKHeightAnchorsakTopakRight Caption   &Bläddra...TabOrderOnClickPuttyPathBrowseButtonClick  	TCheckBoxTelnetForFtpInPuttyCheckLeftToplWidthaHeightAnchorsakLeftakTopakRight Caption2   Öppna &Telnetsessioner i PuTTY för FTP-sessionerTabOrder  TStaticTextPuttyPathHintTextLeft� Top=WidthOHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	   &mönsterTabOrderTabStop	  THistoryComboBoxPuttyRegistryStorageKeyEditLeftTop� WidthjHeightStylecsDropDownListAnchorsakLeftakTopakRight TabOrderOnChangeControlChange    	TTabSheetNetworkSheetTagHelpType	htKeywordHelpKeywordui_pref_networkCaption   Nätverk
ImageIndex
TabVisible
DesignSize��  	TGroupBoxExternalIpAddressGroupBoxLeftTopWidth�HeightbAnchorsakLeftakTopakRight CaptionExtern IP-adressTabOrder 
DesignSize�b  TRadioButtonRetrieveExternalIpAddressButtonLeftTopWidthiHeightAnchorsakLeftakTopakRight Caption/   Hämta extern IP-adress från &operativsystemetTabOrder OnClickControlChange  TRadioButtonCustomExternalIpAddressButtonLeftTop-WidthiHeightAnchorsakLeftakTopakRight Caption%   Använd &följande externa IP-adress:TabOrderOnClickControlChange  TEditCustomExternalIpAddressEditLeft-TopCWidth� HeightTabOrderOnClickControlChange   	TGroupBoxConnectionsGroupLeftToppWidth�Height5AnchorsakLeftakTopakRight CaptionAnslutningarTabOrder
DesignSize�5  	TCheckBoxTryFtpWhenSshFailsCheckLeftTopWidthiHeightAnchorsakLeftakTopakRight Caption-   När SFTP-anslutning av&visas, portknacka FTPTabOrder OnClickControlChange    	TTabSheetPanelRemoteSheetTagHelpType	htKeywordHelpKeywordui_pref_panels_remoteCaption   Fjärr
ImageIndex
TabVisible
DesignSize��  	TGroupBoxPanelsRemoteDirectoryGroupLeftTopWidth�HeightcAnchorsakLeftakTopakRight Caption   FjärrpanelTabOrder 
DesignSize�c  TLabelRefreshRemoteDirectoryUnitLabelLeftPTopEWidthHeightCaptions  	TCheckBoxShowInaccesibleDirectoriesCheckLeftTopWidtheHeightAnchorsakLeftakTopakRight Caption   Vis&a oåtkomliga katalogerTabOrder OnClickControlChange  	TCheckBoxAutoReadDirectoryAfterOpCheckLeftTop-WidtheHeightAnchorsakLeftakTopakRight Caption:Uppdatera auto&matisk katalog efter operation (CTRL+ALT+R)TabOrderOnClickControlChange  	TCheckBoxRefreshRemotePanelCheckLeftTopEWidth
HeightAnchorsakLeftakTopakRight Caption   Uppdatera fjärrpanel varj&eTabOrderOnClickControlChange  TUpDownEditRefreshRemotePanelIntervalEditLeft TopCWidthKHeight	AlignmenttaRightJustify	Increment       �@MaxValue      <�@	MaxLengthTabOrderOnChangeControlChange    	TTabSheetPanelLocalSheetTagHelpType	htKeywordHelpKeywordui_pref_panels_localCaptionLokal
ImageIndex
TabVisible
DesignSize��  	TGroupBoxLocalPanelGroupLeftTopWidth�HeightKAnchorsakLeftakTopakRight CaptionLokal panelTabOrder 
DesignSize�K  	TCheckBoxPreserveLocalDirectoryCheckLeftTopWidtheHeightAnchorsakLeftakTopakRight Caption/   &Ändra inte tillstånd när du byter sessionerTabOrder OnClickControlChange  	TCheckBoxSystemContextMenuCheckLeftTop,WidtheHeightAnchorsakLeftakTopakRight Caption   Använd filsystemets snabbmenyTabOrderOnClickControlChange    	TTabSheetLanguagesSheetTagCaption   Språk
ImageIndex
TabVisible
DesignSize��  	TGroupBoxLanguagesGroupLeftTopWidth�HeightvAnchorsakLeftakTopakRightakBottom Caption   SpråkTabOrder 
DesignSize�v  TLabelLanguageChangeLabelLeftTopXWidth� HeightAnchorsakLeftakBottom Caption-   Ändringar börjar gälla efter nästa start.  	TListViewLanguagesViewLeftTopWidthdHeight5AnchorsakLeftakTopakRightakBottom ColumnsAutoSize	  DoubleBuffered	HideSelectionReadOnly		RowSelect	ParentDoubleBufferedShowColumnHeadersTabOrder 	ViewStylevsReportOnSelectItemListViewSelectItem  TButtonLanguagesGetMoreButtonLeftTopSWidthdHeightAnchorsakRightakBottom Caption   Hämta &fler...TabOrderOnClickLanguagesGetMoreButtonClick     TPanel	LeftPanelLeft Top Width� Height�AlignalLeft
BevelOuterbvNoneTabOrder 
DesignSize� �  	TTreeViewNavigationTreeLeftTop	WidthtHeight�AnchorsakLeftakTopakRightakBottom DoubleBuffered	HideSelectionHotTrack	IndentParentDoubleBufferedReadOnly	ShowButtonsShowRootTabOrder OnChangeNavigationTreeChange
OnChangingNavigationTreeChangingOnCollapsingNavigationTreeCollapsingItems.NodeData
y     6          ��������           E n v i r o n m e n t X 2          ��������            
I n t e r f a c e X ,          ��������            W i n d o w X 2          ��������            
C o m m a n d e r X 0          ��������            	E x p l o r e r X 2          ��������            
L a n g u a g e s X ,          ��������           P a n e l s X ,          ��������            R e m o t e X *          ��������            L o c a l X ,          ��������            E d i t o r X 0          ��������           	T r a n s f e r X 0          ��������            	D r a g D r o p X 4          ��������            B a c k g r o u n d X ,          ��������            R e s u m e X .          ��������            N e t w o r k X 0          ��������            	S e c u r i t y X .          ��������            L o g g i n g X 6       	   ��������           I n t e g r a t i o n X 8          ��������            A p p l i c a t i o n s X 0       
   ��������            	C o m m a n d s X .          ��������            S t o r a g e X .          ��������            U p d a t e s X     TButton
HelpButtonLeft�Top�WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  
TPopupMenuRegisterAsUrlHandlerMenuLeft8Top� 	TMenuItemRegisterAsUrlHandlerItemCaption
RegistreraOnClickRegisterAsUrlHandlerItemClick  	TMenuItemMakeDefaultHandlerItemCaption   Gör WinSCP &standardprogram...OnClickMakeDefaultHandlerItemClick  	TMenuItem!UnregisterForDefaultProtocolsItemCaptionAvregistreraOnClick&UnregisterForDefaultProtocolsItemClick      TPF0TProgressFormProgressFormLeft�Top#HelpType	htKeywordHelpKeywordui_progressBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption	OperationClientHeight� ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnHideFormHideOnShowFormShow
DesignSize��  PixelsPerInch`
TextHeight TLabelOnceDoneOperationLabelLeftBTopXWidthEHeightCaption   När &färdig:FocusControlOnceDoneOperationCombo  TAnimateAnimateLeft
TopWidth-Height<AnchorsakLeftakTopakRight AutoSize	StopFrame  TButtonCancelButtonLeft@TopWidthPHeightAnchorsakTopakRight Cancel	CaptionAvbrytTabOrder OnClickCancelButtonClick  TButtonMinimizeButtonLeft@Top(WidthPHeightAnchorsakTopakRight Caption	&MinimeraTabOrderOnClickMinimizeButtonClick  TPanel	MainPanelLeft
TopAWidth-HeightDAnchorsakLeftakTopakRight 
BevelOuterbvNoneTabOrder
DesignSize-D  TLabelLabel1Left TopWidthHeightCaptionFil:  
TPathLabel	FileLabelLeft8TopWidth� HeightIndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TLabelTargetLabelLeft TopWidth$HeightCaption   Mål:  
TPathLabelTargetPathLabelLeft8TopWidth� HeightIndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TProgressBarTopProgressLeft Top*Width-HeightAnchorsakLeftakTopakRight ParentShowHintShowHint	TabOrder    TPanelTransferPanelLeft
Top� Width-Height?AnchorsakLeftakTopakRight 
BevelOuterbvNoneTabOrder
DesignSize-?  TLabelStartTimeLabelLeftXTopWidthAHeight	AlignmenttaRightJustifyAutoSizeCaption00:00:00  TLabelTimeLeftLabelLeftXTopWidthAHeight	AlignmenttaRightJustifyAutoSizeCaption00:00:00  TLabelTimeLeftLabelLabelLeft TopWidth-HeightCaption	Tid kvar:  TLabelCPSLabelLeft� TopWidthAHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption0 KiB/s  TLabelTimeElapsedLabelLeft� TopWidthAHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption00:00:00  TLabelBytesTransferedLabelLeftXTopWidthAHeight	AlignmenttaRightJustifyAutoSizeCaption0 KiB  TLabelLabel3Left� TopWidthBHeightAnchorsakTopakRight Caption   Förfluten tid:  TLabelStartTimeLabelLabelLeft TopWidth3HeightCaption
Start tid:  TLabelLabel4Left TopWidthYHeightCaption   Bytes överförda:  TLabelLabel12Left� TopWidth"HeightAnchorsakTopakRight Caption
Hastighet:  TProgressBarBottomProgressLeft Top%Width-HeightAnchorsakLeftakTopakRight ParentShowHintShowHint	TabOrder    TPanel
SpeedPanelLeft:Top� Width\Height)AnchorsakTopakRight 
BevelOuterbvNoneTabOrder TLabelSpeedLabel2LeftTop WidthDHeightCaption&Hastighet (kB/s)FocusControl
SpeedCombo  THistoryComboBox
SpeedComboLeftTopWidthPHeightAutoCompleteTabOrder Text
SpeedComboOnExitSpeedComboExit
OnKeyPressSpeedComboKeyPressOnSelectSpeedComboSelectItems.Strings	Unlimited10245122561286432168    	TComboBoxOnceDoneOperationComboLeft@TophWidthPHeightAutoCompleteStylecsDropDownListTabOrder	OnCloseUpOnceDoneOperationComboCloseUpOnSelectOnceDoneOperationComboSelectItems.Strings   Förbli idle   Koppla ifrån   Stäng av dator   TTimerUpdateTimerEnabledOnTimerUpdateTimerTimerLeftPTop�       TPF0TPropertiesDialogPropertiesDialogLeft�Top� HelpType	htKeywordHelpKeywordui_propertiesBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption
PropertiesClientHeight�ClientWidtheColor	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSizee� PixelsPerInch`
TextHeight TButtonOkButtonLeftcTop�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TPageControlPageControlLeftTopWidthZHeightv
ActivePageCommonSheetAnchorsakLeftakTopakRightakBottom TabOrder OnChangePageControlChange 	TTabSheetCommonSheetCaption   Allmänt
DesignSizeRZ  TImageFilesIconImageLeftTopWidth Height Picture.Data
�  TBitmapv  BMv      v   (                    �  �          ��� ��� �� ���  Ɓ  �   w  T  N�  �  w                 3           3333""""""""""3333DDDDDDDDDB 333DDDDDDDDDB333DDDDDDDDDB 33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDDDDB33DDDDDDD  33DDDDDDDBB33DDDDDDD!  33DDDDDDDBB33DDDDDDD!  33DDDDDDDB333!3333DDDDDDD33333333333DDDDDDD33333333333Transparent	  TBevelBevel1LeftTop/Width@Height	AnchorsakLeftakTopakRight Shape	bsTopLine  TLabelLabel1LeftTop:Width,HeightCaptionPlats:  
TPathLabelLocationLabelLeftUTop:Width� HeightUnixPath	IndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TLabel	FileLabelLeftUTopWidth� HeightAutoSizeCaption	FileLabel  TLabelLabel2LeftTopPWidthHeightCaptionStorlek:  TLabel	SizeLabelLeftUTopPWidth� HeightAnchorsakLeftakTopakRight AutoSizeCaption	SizeLabel  TLabelLinksToLabelLabelLeftTopfWidth(HeightCaption   Länkar till:  
TPathLabelLinksToLabelLeftXTopfWidth� HeightUnixPath	IndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TBevelBevel2LeftTop}Width@Height	AnchorsakLeftakTopakRight Shape	bsTopLine  TLabelLabel3LeftTop� Width;HeightCaption   Filrättigheter:FocusControlRightsFrame  TBevelBevel3LeftTop� Width@Height	AnchorsakLeftakTopakRight Shape	bsTopLine  TLabelLabel4LeftTop� Width!HeightCaptionGrupp:FocusControlGroupComboBox  TLabelLabel5LeftTop� Width$HeightCaption   Ägare:FocusControlOwnerComboBox  TImageFileIconImageLeftTopWidth Height   TBevelRecursiveBevelLeftTop8Width@Height	AnchorsakLeftakTopakRight Shape	bsTopLine  �TRightsExtFrameRightsFrameLeftTTop� Width� HeightmTabOrder  	TComboBoxGroupComboBoxLeftUTop� Width� HeightDropDownCount	MaxLength2TabOrderTextGroupComboBoxOnChangeControlChangeOnExitGroupComboBoxExit  	TComboBoxOwnerComboBoxLeftUTop� Width� HeightDropDownCount	MaxLength2TabOrderTextOwnerComboBoxOnChangeControlChangeOnExitOwnerComboBoxExit  	TCheckBoxRecursiveCheckLeftTopBWidth=HeightAnchorsakLeftakTopakRight Caption2   Sätt grupp, ägare och filrättigheter &rekursivtTabOrderOnClickControlChange  TButtonCalculateSizeButtonLeft� TopHWidthPHeightAnchorsakTopakRight Caption	   B&eräknaTabOrder OnClickCalculateSizeButtonClick   	TTabSheetChecksumSheetCaptionKontrollsumma
ImageIndex
DesignSizeRZ  TLabelLabel6LeftTopWidth1HeightCaption
&Algoritm:FocusControlChecksumAlgEdit  	TListViewChecksumViewLeftTop(WidthFHeight)AnchorsakLeftakTopakRightakBottom ColumnsCaptionFilWidth�	WidthType�  CaptionKontrollsummaWidth�	WidthType�   ColumnClickDoubleBuffered	MultiSelect	ReadOnly		RowSelect	ParentDoubleBuffered	PopupMenuListViewMenuTabOrder	ViewStylevsReportOnContextPopupChecksumViewContextPopup  	TComboBoxChecksumAlgEditLeftPTop	WidthyHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeChecksumAlgEditChangeItems.Stringsmd5sha1sha224sha256sha384sha512crc32   TButtonChecksumButtonLeft� TopWidthzHeightAnchorsakTopakRight Caption   B&eräkna kontrollsummaTabOrderOnClickChecksumButtonClick  	TGroupBoxChecksumGroupLeftTop(WidthFHeight)AnchorsakLeftakRightakBottom CaptionKontrollsummaTabOrder
DesignSizeF)  TEditChecksumEditLeft
TopWidth2HeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFaceReadOnly	TabOrder TextChecksumEdit     TButton
HelpButtonLeftTop�WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  
TPopupMenuListViewMenuLeftTop� 	TMenuItemCopyCaption&KopieraOnClick	CopyClick     TPF0TRemoteTransferDialogRemoteTransferDialogLeft(Top� HelpType	htKeywordHelpKeywordui_duplicateBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionRemoteTransferDialogClientHeight� ClientWidthpColor	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSizep�  PixelsPerInch`
TextHeight 	TGroupBoxSymlinkGroupLeftTopWidth`Height� AnchorsakLeftakTopakRightakBottom TabOrder 
DesignSize`�   TLabelSessionLabelLeft1TopWidthJHeightCaption   Mål&session:FocusControlSessionCombo  TLabelLabel2Left1Top<WidthwHeightCaption   Mål för fjärr&katalog:FocusControlDirectoryEdit  TImageImageLeftTopWidth Height AutoSize	Picture.Data
�  	TPngImage�PNG

   IHDR           szz�   	pHYs  �  ��o�d  mIDATx���LSW��m�ƍ�.f��#�2���dL������ ��s s>X@1�0���1[&n�b�h�����(�l]��C;hזR�����Z)}x[Yv�����|�w�{�wZ
�s�\o[�I��,v$Is⌓(��6��t��ohU5[�$�q ��[".u@7j��^�c#< 67@o���A����4!�j&_	�`�9���ŀ�f�A?j����Ah]�[��<��N(�+�@*DKa�:9�* ��q��=�=��-	�Y�#�ʉ�q́�u?P����
��1��*�՛�� ��Β�a0;8t�OCP���%$�&��Xq�HrW`�dGAݹG߂iO;�ߺ� D卤&o%t4�K�S߄ɪ@��I"�O�����~��>V,�u�'�-Z;)u�d�;Ad����8-��ᥘ����u1c^,'�ĺA���Y�Z7 ��8�~�����J��"9}����Y��on��#*����<�n0��v7ٶ4������%�3 �Ǉ�D�z��#S���R��a~�y�b��R�,��/��ȶ��zԎby��@��|7 � v'��kw�{�)t>��5�U7�T�q��Ϻ� >!����.� ��A(>�
5�o,J9��9������ �,!��>Nj"�}	��3��� :���w|q�r�V쯿i޻,��tIN�O(6�;�W�=��}�΂�sJD,�DTl��/��~�e�) �ë���|�ؾ���n�W�g(
�)p`��ĥ�$P{򭫂��@ ׹�������9X�v�g
kO�n�j_���(��=p��m(n����cb�0�9IO���4 �E���-h���m�kX_^���$�H >\0 �ފVz*���� ���K�rp_�? D^�����1�q{T�t5�����aƳI���K���O���T�|�0;|�ޭ��ӄ_Ht�0F��ﱀ��mIF� ���R�������@0-�s,qu���`6�\��f1:��pҙ�Ҿ�a��UGqtofh -��������b��	�nŕ��~_v�����0#z�֙1!M���a��`���j��{9���B��A�_���[?�nF�    IEND�B`�  	TComboBoxSessionComboLeft1TopWidth$HeightStylecsDropDownListAnchorsakLeftakTopakRight DropDownCount	MaxLength� TabOrder OnChangeSessionComboChange  THistoryComboBoxDirectoryEditLeft1TopLWidth$HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChange  	TCheckBoxNotDirectCopyCheckLeft7TopiWidth HeightAnchorsakLeftakTopakRight Caption"   Dubblera via lokal temporär kopiaTabOrderOnClickNotDirectCopyCheckClick   TButtonOkButtonLefttTop� WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top� WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeftTop� WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick    TPF0�TRightsExtFrameRightsExtFrameWidth� Heightm �TLabel
OctalLabelLeftTopDWidthHeightCaptionO&ktal:FocusControl	OctalEdit  �TGrayedCheckBoxGroupReadCheckTabOrder  �TGrayedCheckBoxGroupWriteCheckTabOrder  �TGrayedCheckBoxGroupExecuteCheckTabOrder  �TGrayedCheckBoxOthersReadCheckTabOrder  �TGrayedCheckBoxOthersWriteCheckTabOrder	  �TGrayedCheckBoxOthersExecuteCheckTabOrder
  �	TCheckBoxDirectoriesXCheckTopYTabOrder  �TEdit	OctalEditLeft7Top@Width@Height	MaxLengthTabOrderText	OctalEditOnChangeOctalEditChangeOnExitOctalEditExit  �TGrayedCheckBoxSetUidCheckTag Left� TopWidthFHeightCaption	   Sätt UIDTabOrderOnClickControlChange  �TGrayedCheckBoxSetGIDCheckTag Left� TopWidthFHeightCaption	   Sätt GIDTabOrderOnClickControlChange  �TGrayedCheckBoxStickyBitCheckTag Left� Top+WidthFHeightCaption
Sticky bitTabOrderOnClickControlChange  �TButtonCloseButtonLeft� TopPWidthKHeightCaption   StängTabOrderVisibleOnClickCloseButtonClick   TPF0TRightsFrameRightsFrameLeft Top Width� HeightWTabOrder OnContextPopupFrameContextPopup TLabel
OwnerLabelLeftTopWidth HeightCaption   &ÄgareFocusControlOwnerReadCheck  TLabel
GroupLabelLeftTopWidthHeightCaption&GruppFocusControlGroupReadCheck  TLabelOthersLabelLeftTop,Width!HeightCaptionA&ndraFocusControlOthersReadCheck  TSpeedButtonOthersButtonTagLeft Top)Width8HeightFlat	OnClickRightsButtonsClick  TSpeedButtonGroupButtonTagLeft TopWidth8HeightFlat	OnClickRightsButtonsClick  TSpeedButtonOwnerButtonTagLeft TopWidth8HeightFlat	OnClickRightsButtonsClick  TGrayedCheckBoxOwnerReadCheckTag Left:TopWidth"HeightHint   LäsCaptionRParentShowHintShowHint	TabOrder OnClickControlChange  TGrayedCheckBoxOwnerWriteCheckTag� Left_TopWidth"HeightHintSkrivCaptionWParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxOwnerExecuteCheckTag@Left� TopWidthHeightHint   Kör/ÖppnaCaptionXParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxGroupReadCheckTag Left:TopWidth"HeightCaptionRParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxGroupWriteCheckTagLeft_TopWidth!HeightCaptionWParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxGroupExecuteCheckTagLeft� TopWidthHeightCaptionXParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxOthersReadCheckTagLeft:Top+Width"HeightCaptionRParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxOthersWriteCheckTagLeft_Top+Width!HeightCaptionWParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxOthersExecuteCheckTagLeft� Top+WidthHeightCaptionXParentShowHintShowHint	TabOrderOnClickControlChange  	TCheckBoxDirectoriesXCheckLeftTopAWidth� HeightCaptionAddera &X till katalogerTabOrder	OnClickControlChange  
TPopupMenuRightsPopupImagesRightsImagesOnPopupRightsPopupPopupLeft� Top; 	TMenuItem	Norights1ActionNoRightsAction  	TMenuItemDefaultrights1ActionDefaultRightsAction  	TMenuItem
Allrights1ActionAllRightsAction  	TMenuItem
Leaveasis1ActionLeaveRightsAsIsAction  	TMenuItemN1Caption-  	TMenuItemCopyAsText1ActionCopyTextAction  	TMenuItemCopyAsOctal1ActionCopyOctalAction  	TMenuItemPaste1ActionPasteAction   TActionListRightsActionsImagesRightsImages	OnExecuteRightsActionsExecuteOnUpdateRightsActionsUpdateLeft� Top TActionNoRightsActionCaption   I&nga rättigheter
ImageIndex ShortCutN@  TActionDefaultRightsActionCaption   Stan&dardrättigheter
ImageIndexShortCutD@  TActionAllRightsActionCaption   &Alla rättigheter
ImageIndexShortCutA@  TActionLeaveRightsAsIsActionCaption   &Lämna oförändradShortCutL@  TActionCopyTextActionCaption&Kopiera som text
ImageIndexShortCutC@  TActionCopyOctalActionCaptionKopiera som &oktalt
ImageIndexShortCutO@  TActionPasteActionCaptionKl&istra in
ImageIndexShortCutV@   TPngImageListRightsImages	PngImages
BackgroundclWindowName'No rights-preset on permissions controlPngImage.Data
l  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�}�mH�Q��ϳ��^ܴ�h�--�1]bm�l}�̂�ä~��b�$AIER �EJ��6ɷ�N�d�/ihkj{s�����`��u�r�=���9��s)l�N���%�@��RI�X�YL{n�L&?��/�����O���慃p ��S5E��;�����"z�X�~Fl�d�4�Մdi��X �N��>��<����.�d�������2�k�pb�e��JU!R��tR�#��P1D�g����x�|~�\��W��4[6�ey��8k�`ܩ��t�G���y�P��asa|��=C�*+�H����},�61c�vY���8�Z��@���+���E�ç���l=������y����;B �G��Tub:�9�eg��X��@A{{�����۶=��C��=��g�d��FU����]x�ܫP�����<l?���>O�:���I8���! ��g���+������r�.]�t~��IX �$��1�u+O}��S��� �%<ilB��8�N���!]&A
	�Y^�m�Y������XƧ8��E�+�H	`<_�����1�r!Y*����}��.�!02a�#�L�C�铈_ZD�(
_<^�E���fʤs��{c�~�F�EKp�(�zd��p0����N�Ǒ��$[�#�Z(�P  
����h=�%�s`�S�v;����7�.��$+��,Ҁ    IEND�B`� 
BackgroundclWindowNameDefault rights-presetPngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  mIDATx�cd����x�����@|��?�Jn�/��R���t����{/�iŀ	�q3~u�� S{�F Uď��K���s������L�br@�t���z���{�J�0108�<�u?L������>��;�nU���̷7\�W������e�����t3V��� �� �Mg���1�J(�?��
�ٸ�33�<,���-���{��e�)f�FV�@��3׈7`�s@MP@:p�2��=z����4?�a��`W�>r�x����0;�aƜ�`��g�7����`M9�	s,�`Ӟ��p��-��a��n�1�8w�.B3ԀU[�7�℄-y� :���    IEND�B`� 
BackgroundclWindowNameAll rights-presetPngImage.Data
@  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڅ�HSQǿ�mӵ7*i�$ڔ�b���A��U��0���!B*�!T&%iEP3�DB0J�B݆��sj�j��GK�ԙn2������H���{�9�s�{�RX�Z-���+��L�� :��dh�-����B��9���I��43���Z������c�xh��a�	E��Y8�q7��ڼ5	*� 적CfcM�3Q�9�$�a1�D���/��s����W�N�"#@"��'&�j��
8�ͱ����!�ڪJ��u�������<]�Õ\�^�o���!
|jn��/������>9;���uu����v��?�������? b7Y{W�������*��\kY�ԙl$i��%�����m�HI�ךu�D�1]25�m�/M#~��$I���u(-�D�|ƾ�`��2&W���HwnW��^o�̤'�`4w�U���1.=φ���ͬ���Ao+FRV"ۆ�g�T�,���4���E�8*�O1D��I��`�3������`y��z�s1���������D#-_q� !���i�wvѪH����hX���Ӆ��F[�g��A�a���(E���a�sc�a��t��Ĉ��u))!ʽr�V� Q
!��Q7�����2�A����z"�n�/��&�<��Y��]�����\UɅ    IEND�B`� 
BackgroundclWindowNameCopy rights-permissions as textPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  IDATxڍ��KSQǿ�%5zQF��A���ڃ= D���>̱��Q�V������Z�(JɈ�ħ��$����L�f�����8E�������p�pB.�>"���+șB5�Y�T��H���)r�����n���"��#y�[T�
8w�	_.E��O݁�l�e�M�Ðo�f���-Iv�a}�Pl4���:�����HG����3�	"���n( ��'t%8Q��I������������"���D�
���B���=}�}���N��`�s8\{$#��;$�������.�������D8|=$�[`碸�:��R�:����g��]������`��&�`��o�5���Ch�h����?�b��ڹJpR��ؐ�nˇ|�$�N��j�:�ZX��q`�:u_9�h���ņ̦$������1�E0�{���[�Dʥ��� 98*����Y� �Хs"��9.����ڇ.����1�Zض��8� �A��i�fv WS�)�_�    IEND�B`� 
BackgroundclWindowName Copy rights-permissions as octalPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?Cf���X�1&���Ӳþ`��e=��(�g���?�����t���VC��w��?�,����(
>}��p��+���/�c`fu�U���i����,b���/X�t�6�>B�܀��5�gU�0|�1�l�b�7 �u���U�^aX����n/�z�<�K3�}ހHj^�Vu8CL�����S62̪�{	xؙ^���p��+���]�]�6 �i���Ց�Us&�$0T�@x	��y�p��S0�νGs*C��7,�?�&�!�zÄ���)���a��f��_b���æ�g�V�A��[�Vm4�ƃ���>����ˀ�%�n�g����n��y�bj�ex��XAݔ5�^���`��9���EA������YX���m�l]޿�aaC4� FFF����]��%t5�{+���2��s0,j��n@t�/aU���4�c7 �j�"���D��   ,E��d�    IEND�B`� 
BackgroundclWindowNamePastePngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�cd@���]�����3L߸qm���	����?�#��]@Cmذ6�3��iǪ|��c�~0扌��-���79��Ǘ���cЛ��p���Ƿ�2 `�j�kx0�ۧ�Q$�}K���cL�ݧe�}��2�	�_f��3���.�(G.?dX���1&�_`C�8�1�ytŀ�ߓf�2|��E�ӗ�W�fX���9fVw�N!���_GQ��g2ì�`��Y�b��<��/�e�r�Ê]箂p�gxq�����a���/���;/�_{
f߹���n_AQ��_*��P�������æ�g ���2<�qE�2�4�Y�����j����m�`������E�Y�fWG2T����Hk����l��]>��`[&��(�w_�0���� H��3|z�Er�x9ì�h�����j.
�b��[����a�z��o��vAU�rF\�QU��3 
+�Ed��    IEND�B`�  Left� Bitmap
        TPF0�TScpCommanderFormScpCommanderFormLeft� Top HelpType	htKeywordHelpKeywordui_commanderCaptionScpCommanderFormClientHeight�ClientWidth=OldCreateOrder	PixelsPerInch`
TextHeight � 	TSplitterSplitterLeft�Top� WidthHeight*CursorcrSizeWEHintj   |Dra för att ändra proportioner på filpaneler. Dubbelklicka för att bredden på filpanelerna ska lika.ResizeStylersUpdateOnCanResizeSplitterCanResizeOnMovedSplitterMoved  �	TSplitterQueueSplitterTopWidth=  �TTBXDockTopDockWidth=Height�  TTBXToolbarMenuToolbarLeft Top CaptionMenyCloseButtonImagesGlyphsModule.ExplorerImagesMenuBar	
ShrinkModetbsmWrapStretch	TabOrder TTBXSubmenuItemLocalMenuButtonCaption&LokalHelpKeywordui_commander_menu#localHintC   Ändra layout för lokal panel eller ändra katalog/enhet som visas TTBXItemTBXItem1Action)NonVisualDataModule.LocalChangePathAction  TTBXSeparatorItemTBXSeparatorItem1  TTBXSubmenuItemTBXSubmenuItem2Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItemTBXItem2Action&NonVisualDataModule.LocalOpenDirAction  TTBXItemTBXItem3Action/NonVisualDataModule.LocalExploreDirectoryAction  TTBXSeparatorItemTBXSeparatorItem2  TTBXItemTBXItem4Action(NonVisualDataModule.LocalParentDirAction  TTBXItemTBXItem5Action&NonVisualDataModule.LocalRootDirAction  TTBXItemTBXItem6Action&NonVisualDataModule.LocalHomeDirAction  TTBXSeparatorItemTBXSeparatorItem3  TTBXItemTBXItem7Action#NonVisualDataModule.LocalBackAction  TTBXItemTBXItem8Action&NonVisualDataModule.LocalForwardAction   TTBXItemTBXItem9Action&NonVisualDataModule.LocalRefreshAction  TTBXItem	TBXItem10Action*NonVisualDataModule.LocalAddBookmarkAction  TTBXItem	TBXItem11Action.NonVisualDataModule.LocalPathToClipboardAction  TTBXSeparatorItemTBXSeparatorItem4  TTBXSubmenuItemTBXSubmenuItem3Caption&SorteraHelpKeywordui_file_panel#sorting_filesHint   Ändra filordning i lokal panel TTBXItem	TBXItem12Action,NonVisualDataModule.LocalSortAscendingAction  TTBXSeparatorItemTBXSeparatorItem5  TTBXItem	TBXItem13Action)NonVisualDataModule.LocalSortByNameAction
GroupIndex	RadioItem	  TTBXItem	TBXItem14Action(NonVisualDataModule.LocalSortByExtAction
GroupIndex	RadioItem	  TTBXItem	TBXItem15Action)NonVisualDataModule.LocalSortByTypeAction
GroupIndex	RadioItem	  TTBXItem	TBXItem16Action,NonVisualDataModule.LocalSortByChangedAction
GroupIndex	RadioItem	  TTBXItem	TBXItem17Action)NonVisualDataModule.LocalSortBySizeAction
GroupIndex	RadioItem	  TTBXItem	TBXItem18Action)NonVisualDataModule.LocalSortByAttrAction
GroupIndex	RadioItem	   TTBXSubmenuItemTBXSubmenuItem4Caption&Visa kolumnerHelpKeywordui_file_panel#selecting_columnsHint$   Välj kolumner som ska visas i panel TTBXItem	TBXItem19Action1NonVisualDataModule.ShowHideLocalNameColumnAction  TTBXItem	TBXItem20Action1NonVisualDataModule.ShowHideLocalSizeColumnAction  TTBXItem	TBXItem21Action1NonVisualDataModule.ShowHideLocalTypeColumnAction  TTBXItem	TBXItem22Action4NonVisualDataModule.ShowHideLocalChangedColumnAction  TTBXItem	TBXItem23Action1NonVisualDataModule.ShowHideLocalAttrColumnAction   TTBXItem
TBXItem221Action%NonVisualDataModule.LocalFilterAction   TTBXSubmenuItemTBXSubmenuItem18Caption&MarkeraHelpKeywordui_commander_menu#markHint   Kommandon för markera TTBXItem
TBXItem107Action#NonVisualDataModule.SelectOneAction  TTBXItem
TBXItem108Action NonVisualDataModule.SelectAction  TTBXItem
TBXItem109Action"NonVisualDataModule.UnselectAction  TTBXItem
TBXItem110Action#NonVisualDataModule.SelectAllAction  TTBXItem
TBXItem111Action)NonVisualDataModule.InvertSelectionAction  TTBXItem
TBXItem112Action(NonVisualDataModule.ClearSelectionAction  TTBXItem	TBXItem27Action*NonVisualDataModule.RestoreSelectionAction   TTBXSubmenuItemTBXSubmenuItem5Caption&FilerHelpKeywordui_commander_menu#filesHint   Kommandon för filoperationer TTBXSubmenuItemTBXSubmenuItem26Caption&NyHelpKeyword
task_indexHintSkapa objekt|Skapa nytt objekt TTBXItem	TBXItem28Action!NonVisualDataModule.NewFileAction  TTBXItem	TBXItem24Action NonVisualDataModule.NewDirAction  TTBXItem
TBXItem209Action!NonVisualDataModule.NewLinkAction   TTBXSeparatorItemTBXSeparatorItem6  TTBXItem	TBXItem25Action%NonVisualDataModule.CurrentOpenAction  TTBXItem	TBXItem26Action%NonVisualDataModule.CurrentEditAction  TTBXSubmenuItemTBXSubmenuItem25Action0NonVisualDataModule.CurrentEditAlternativeAction  TTBXItem	TBXItem29Action,NonVisualDataModule.CurrentAddEditLinkAction  TTBXSeparatorItemTBXSeparatorItem7  TTBXItemCurrentCopyItemAction$NonVisualDataModule.RemoteCopyAction  TTBXItemCurrentMoveItemAction$NonVisualDataModule.RemoteMoveAction  TTBXItem	TBXItem31Action&NonVisualDataModule.RemoteCopyToAction  TTBXItem	TBXItem33Action&NonVisualDataModule.RemoteMoveToAction  TTBXItem	TBXItem34Action'NonVisualDataModule.CurrentDeleteAction  TTBXItem	TBXItem35Action'NonVisualDataModule.CurrentRenameAction  TTBXItem	TBXItem36ActionNonVisualDataModule.PasteAction  TTBXSeparatorItemTBXSeparatorItem8  TTBXSubmenuItemCustomCommandsMenuAction(NonVisualDataModule.CustomCommandsAction  TTBXSubmenuItemTBXSubmenuItem6Caption&FilnamnHelpKeyword	filenamesHint$   Operationer med namn på valda filer TTBXItem	TBXItem37Action/NonVisualDataModule.FileListToCommandLineAction  TTBXItem	TBXItem38Action-NonVisualDataModule.FileListToClipboardAction  TTBXItem	TBXItem39Action1NonVisualDataModule.FullFileListToClipboardAction  TTBXItem	TBXItem40Action(NonVisualDataModule.UrlToClipboardAction   TTBXSeparatorItemTBXSeparatorItem9  TTBXItem	TBXItem41Action+NonVisualDataModule.CurrentPropertiesAction   TTBXSubmenuItemTBXSubmenuItem7Caption
&KommandonHelpKeywordui_commander_menu#commandsHintAndra kommandon TTBXItem	TBXItem42Action,NonVisualDataModule.CompareDirectoriesAction  TTBXItem	TBXItem43Action%NonVisualDataModule.SynchronizeAction  TTBXItem	TBXItem44Action)NonVisualDataModule.FullSynchronizeAction  TTBXItem	TBXItem45Action-NonVisualDataModule.SynchronizeBrowsingAction  TTBXItem
TBXItem210Action)NonVisualDataModule.RemoteFindFilesAction  TTBXSubmenuItemQueueSubmenuItemCaption   K&öHelpKeywordui_queue#managing_the_queueHint   Kommandon för kölistaOnPopupQueueSubmenuItemPopup TTBXItemQueueEnableItem2Action%NonVisualDataModule.QueueEnableAction  TTBXItem	TBXItem46Action#NonVisualDataModule.QueueGoToAction  TTBXSeparatorItemTBXSeparatorItem10  TTBXItem	TBXItem47Action(NonVisualDataModule.QueueItemQueryAction  TTBXItem	TBXItem48Action(NonVisualDataModule.QueueItemErrorAction  TTBXItem	TBXItem49Action)NonVisualDataModule.QueueItemPromptAction  TTBXSeparatorItemTBXSeparatorItem11  TTBXItem	TBXItem50Action*NonVisualDataModule.QueueItemExecuteAction  TTBXItem
TBXItem196Action(NonVisualDataModule.QueueItemPauseAction  TTBXItem
TBXItem197Action)NonVisualDataModule.QueueItemResumeAction  TTBXItem	TBXItem51Action)NonVisualDataModule.QueueItemDeleteAction  TTBXComboBoxItemQueueSpeedComboBoxItemAction(NonVisualDataModule.QueueItemSpeedAction  TTBXSeparatorItemTBXSeparatorItem12  TTBXItem	TBXItem52Action%NonVisualDataModule.QueueItemUpAction  TTBXItem	TBXItem53Action'NonVisualDataModule.QueueItemDownAction  TTBXSeparatorItemTBXSeparatorItem48  TTBXSubmenuItemTBXSubmenuItem13Caption&AllaHelpKeywordui_queue#managing_the_queueHint&   Administrationskommandon för kömassa TTBXItem
TBXItem198Action'NonVisualDataModule.QueuePauseAllAction  TTBXItem
TBXItem199Action(NonVisualDataModule.QueueResumeAllAction  TTBXSeparatorItemTBXSeparatorItem39  TTBXItem
TBXItem134Action,NonVisualDataModule.QueueDeleteAllDoneAction    TTBXSeparatorItemTBXSeparatorItem13  TTBXItem	TBXItem54Action!NonVisualDataModule.ConsoleAction  TTBXItem	TBXItem55ActionNonVisualDataModule.PuttyAction  TTBXSeparatorItemTBXSeparatorItem14  TTBXItem	TBXItem56Action(NonVisualDataModule.FileSystemInfoAction  TTBXItem	TBXItem57Action%NonVisualDataModule.ClearCachesAction  TTBXSeparatorItemTBXSeparatorItem15  TTBXItem	TBXItem58Action*NonVisualDataModule.CloseApplicationAction   TTBXSubmenuItemTBXSubmenuItem19Caption&SessionHelpKeywordui_commander_menu#sessionHint   Kommandon för session TTBXItem
TBXItem113Action$NonVisualDataModule.NewSessionAction  TTBXItem
TBXItem218Action*NonVisualDataModule.DuplicateSessionAction  TTBXItem
TBXItem115Action&NonVisualDataModule.CloseSessionAction  TTBXItem
TBXItem114Action-NonVisualDataModule.SaveCurrentSessionAction2  TTBXSeparatorItemTBXSeparatorItem29  TTBXSubmenuItemTBXSubmenuItem21Action(NonVisualDataModule.OpenedSessionsAction  TTBXSubmenuItemTBXSubmenuItem231Action$NonVisualDataModule.WorkspacesAction  TTBXItem
TBXItem230Action'NonVisualDataModule.SaveWorkspaceAction  TTBXSeparatorItemTBXSeparatorItem53  TTBXSubmenuItemTBXSubmenuItem20Action(NonVisualDataModule.SavedSessionsAction2   TTBXSubmenuItemTBXSubmenuItem9Caption&AlternativHelpKeywordui_commander_menu#optionsHint)   Ändra layout/inställningar för program TTBXSubmenuItemTBXSubmenuItem10Caption   &VerktygsfältHelpKeywordui_toolbarsHint   Visa/dölj verktygsfält TTBXItem	TBXItem64Action/NonVisualDataModule.CommanderCommandsBandAction  TTBXItem	TBXItem60Action.NonVisualDataModule.CommanderSessionBandAction  TTBXItem	TBXItem62Action2NonVisualDataModule.CommanderPreferencesBandAction  TTBXItem	TBXItem63Action+NonVisualDataModule.CommanderSortBandAction  TTBXItem
TBXItem186Action.NonVisualDataModule.CommanderUpdatesBandAction  TTBXItem
TBXItem188Action/NonVisualDataModule.CommanderTransferBandAction  TTBXItem
TBXItem215Action5NonVisualDataModule.CommanderCustomCommandsBandAction  TTBXSeparatorItemTBXSeparatorItem38  TTBXItem	TBXItem74Action"NonVisualDataModule.ToolBar2Action  TTBXSeparatorItemTBXSeparatorItem47  TTBXItem
TBXItem191Action&NonVisualDataModule.LockToolbarsAction  TTBXItem
TBXItem133Action.NonVisualDataModule.SelectiveToolbarTextAction   TTBXSubmenuItemTBXSubmenuItem11Caption&Lokal panelHelpKeywordui_file_panelHint   Ändra layout för lokal panel TTBXItem	TBXItem65Action3NonVisualDataModule.CommanderLocalHistoryBandAction  TTBXItem	TBXItem66Action6NonVisualDataModule.CommanderLocalNavigationBandAction  TTBXItem	TBXItem59Action0NonVisualDataModule.CommanderLocalFileBandAction  TTBXItem	TBXItem61Action5NonVisualDataModule.CommanderLocalSelectionBandAction  TTBXSeparatorItemTBXSeparatorItem16  TTBXItem	TBXItem67Action#NonVisualDataModule.LocalTreeAction  TTBXSeparatorItemTBXSeparatorItem17  TTBXItem	TBXItem68Action(NonVisualDataModule.LocalStatusBarAction   TTBXSubmenuItemTBXSubmenuItem12Caption   F&järrpanelHelpKeywordui_file_panelHint   Ändra layout för fjärrpanel TTBXItem	TBXItem69Action4NonVisualDataModule.CommanderRemoteHistoryBandAction  TTBXItem	TBXItem70Action7NonVisualDataModule.CommanderRemoteNavigationBandAction  TTBXItem
TBXItem136Action1NonVisualDataModule.CommanderRemoteFileBandAction  TTBXItem
TBXItem131Action6NonVisualDataModule.CommanderRemoteSelectionBandAction  TTBXSeparatorItemTBXSeparatorItem18  TTBXItem	TBXItem71Action$NonVisualDataModule.RemoteTreeAction  TTBXSeparatorItemTBXSeparatorItem19  TTBXItem	TBXItem72Action)NonVisualDataModule.RemoteStatusBarAction   TTBXSeparatorItemTBXSeparatorItem20  TTBXItemSessionsTabsAction3Action&NonVisualDataModule.SessionsTabsAction  TTBXItem	TBXItem73Action*NonVisualDataModule.CommandLinePanelAction  TTBXItem	TBXItem75Action#NonVisualDataModule.StatusBarAction  TTBXItem	TBXItem76Action!NonVisualDataModule.ViewLogAction  TTBXSubmenuItemTBXSubmenuItem14Caption   K&öHelpKeywordui_queueHint   Konfigurera kölista TTBXItem	TBXItem77Action#NonVisualDataModule.QueueShowAction	RadioItem	  TTBXItem	TBXItem78Action,NonVisualDataModule.QueueHideWhenEmptyAction	RadioItem	  TTBXItem	TBXItem79Action#NonVisualDataModule.QueueHideAction	RadioItem	  TTBXSeparatorItemTBXSeparatorItem21  TTBXItem	TBXItem80Action&NonVisualDataModule.QueueToolbarAction  TTBXSeparatorItemTBXSeparatorItem22  TTBXSubmenuItemTBXSubmenuItem8Action-NonVisualDataModule.QueueCycleOnceEmptyActionDropdownCombo	 TTBXItem
TBXItem222Action,NonVisualDataModule.QueueIdleOnceEmptyAction	RadioItem	  TTBXItem
TBXItem223Action2NonVisualDataModule.QueueDisconnectOnceEmptyAction	RadioItem	  TTBXItem
TBXItem224Action0NonVisualDataModule.QueueShutDownOnceEmptyAction	RadioItem	   TTBXItem	TBXItem81Action*NonVisualDataModule.QueuePreferencesAction   TTBXSeparatorItemTBXSeparatorItem23  TTBXColorItemColorMenuItemAction#NonVisualDataModule.ColorMenuActionColorclNone  TTBXSeparatorItemTBXSeparatorItem49  TTBXItem	TBXItem82Action%NonVisualDataModule.PreferencesAction   TTBXSubmenuItemRemoteMenuButtonCaption   F&järrHelpKeywordui_commander_menu#remoteHint=   Ändra layout för fjärrpanel eller ändra katalog som visas TTBXItem	TBXItem83Action*NonVisualDataModule.RemoteChangePathAction  TTBXSeparatorItemTBXSeparatorItem24  TTBXSubmenuItemTBXSubmenuItem15Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItem	TBXItem84Action'NonVisualDataModule.RemoteOpenDirAction  TTBXSeparatorItemTBXSeparatorItem25  TTBXItem	TBXItem85Action)NonVisualDataModule.RemoteParentDirAction  TTBXItem	TBXItem86Action'NonVisualDataModule.RemoteRootDirAction  TTBXItem	TBXItem87Action'NonVisualDataModule.RemoteHomeDirAction  TTBXSeparatorItemTBXSeparatorItem26  TTBXItem	TBXItem88Action$NonVisualDataModule.RemoteBackAction  TTBXItem	TBXItem89Action'NonVisualDataModule.RemoteForwardAction   TTBXItem	TBXItem90Action'NonVisualDataModule.RemoteRefreshAction  TTBXItem	TBXItem91Action+NonVisualDataModule.RemoteAddBookmarkAction  TTBXItem	TBXItem92Action/NonVisualDataModule.RemotePathToClipboardAction  TTBXSeparatorItemTBXSeparatorItem27  TTBXSubmenuItemTBXSubmenuItem16Caption&SorteraHelpKeywordui_file_panel#sorting_filesHint   Ändra filordning i fjärrpanel TTBXItem	TBXItem93Action-NonVisualDataModule.RemoteSortAscendingAction  TTBXSeparatorItemTBXSeparatorItem28  TTBXItem	TBXItem94Action*NonVisualDataModule.RemoteSortByNameAction
GroupIndex	RadioItem	  TTBXItem	TBXItem95Action)NonVisualDataModule.RemoteSortByExtAction
GroupIndex	RadioItem	  TTBXItem
TBXItem193Action*NonVisualDataModule.RemoteSortByTypeAction	RadioItem	  TTBXItem	TBXItem96Action-NonVisualDataModule.RemoteSortByChangedAction
GroupIndex	RadioItem	  TTBXItem	TBXItem97Action*NonVisualDataModule.RemoteSortBySizeAction
GroupIndex	RadioItem	  TTBXItem	TBXItem98Action,NonVisualDataModule.RemoteSortByRightsAction
GroupIndex	RadioItem	  TTBXItem	TBXItem99Action+NonVisualDataModule.RemoteSortByOwnerAction
GroupIndex	RadioItem	  TTBXItem
TBXItem100Action+NonVisualDataModule.RemoteSortByGroupAction
GroupIndex	RadioItem	   TTBXSubmenuItemTBXSubmenuItem17Caption&Visa kolumnerHelpKeywordui_file_panel#selecting_columnsHint$   Välj kolumner som ska visas i panel TTBXItem
TBXItem101Action2NonVisualDataModule.ShowHideRemoteNameColumnAction  TTBXItem
TBXItem102Action2NonVisualDataModule.ShowHideRemoteSizeColumnAction  TTBXItem
TBXItem192Action2NonVisualDataModule.ShowHideRemoteTypeColumnAction  TTBXItem
TBXItem103Action5NonVisualDataModule.ShowHideRemoteChangedColumnAction  TTBXItem
TBXItem104Action4NonVisualDataModule.ShowHideRemoteRightsColumnAction  TTBXItem
TBXItem105Action3NonVisualDataModule.ShowHideRemoteOwnerColumnAction  TTBXItem
TBXItem106Action3NonVisualDataModule.ShowHideRemoteGroupColumnAction  TTBXItem
TBXItem179Action8NonVisualDataModule.ShowHideRemoteLinkTargetColumnAction   TTBXItem
TBXItem220Action&NonVisualDataModule.RemoteFilterAction   TTBXSubmenuItemTBXSubmenuItem22Caption   &HjälpHelpKeywordui_commander_menu#helpHint   Hjälp TTBXItem
TBXItem116Action)NonVisualDataModule.TableOfContentsAction  TTBXSeparatorItemTBXSeparatorItem30  TTBXItem
TBXItem117Action"NonVisualDataModule.HomepageAction  TTBXItem
TBXItem118Action#NonVisualDataModule.ForumPageAction  TTBXItem
TBXItem119Action%NonVisualDataModule.HistoryPageAction  TTBXSeparatorItemTBXSeparatorItem31  TTBXItem
TBXItem120Action)NonVisualDataModule.CheckForUpdatesAction  TTBXSeparatorItemTBXSeparatorItem32  TTBXItem
TBXItem121Action$NonVisualDataModule.DonatePageAction  TTBXSeparatorItemTBXSeparatorItem33  TTBXItem
TBXItem122ActionNonVisualDataModule.AboutAction    TTBXToolbarPreferencesToolbarLeft Top3Caption   InställningarDockPos DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem126Action%NonVisualDataModule.PreferencesAction  TTBXSeparatorItemTBXSeparatorItem36  TTBXItem
TBXItem127Action!NonVisualDataModule.ViewLogAction  TTBXSubmenuItemTBXSubmenuItem24Action)NonVisualDataModule.QueueToggleShowActionDisplayModenbdmImageAndTextDropdownCombo	 TTBXItem
TBXItem128Action#NonVisualDataModule.QueueShowAction	RadioItem	  TTBXItem
TBXItem129Action,NonVisualDataModule.QueueHideWhenEmptyAction	RadioItem	  TTBXItem
TBXItem130Action#NonVisualDataModule.QueueHideAction	RadioItem	    TTBXToolbarSessionToolbarLeft TopCaptionSessionDockPos DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder  TTBXItem
TBXItem123Action$NonVisualDataModule.NewSessionActionDisplayModenbdmImageAndText  TTBXItem
TBXItem219Action*NonVisualDataModule.DuplicateSessionAction  TTBXItem
TBXItem124Action&NonVisualDataModule.CloseSessionAction  TTBXItem
TBXItem125Action-NonVisualDataModule.SaveCurrentSessionAction2  TTBXSeparatorItemTBXSeparatorItem34  TTBXSubmenuItemTBXSubmenuItem23Action(NonVisualDataModule.SavedSessionsAction2DisplayModenbdmImageAndTextOptionstboDropdownArrow    TTBXToolbarSortToolbarLeft TopMCaptionSorteraDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem145Action.NonVisualDataModule.CurrentSortAscendingAction  TTBXSeparatorItemTBXSeparatorItem40  TTBXItem
TBXItem146Action+NonVisualDataModule.CurrentSortByNameAction  TTBXItem
TBXItem147Action*NonVisualDataModule.CurrentSortByExtAction  TTBXItem
TBXItem148Action+NonVisualDataModule.CurrentSortByTypeAction  TTBXItem
TBXItem149Action.NonVisualDataModule.CurrentSortByChangedAction  TTBXItem
TBXItem150Action+NonVisualDataModule.CurrentSortBySizeAction  TTBXItem
TBXItem151Action-NonVisualDataModule.CurrentSortByRightsAction  TTBXItem
TBXItem152Action,NonVisualDataModule.CurrentSortByOwnerAction  TTBXItem
TBXItem153Action,NonVisualDataModule.CurrentSortByGroupAction   TTBXToolbarCommandsToolbarLeft TopgCaption	KommandonDockPos DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem154Action,NonVisualDataModule.CompareDirectoriesAction  TTBXItem
TBXItem155Action%NonVisualDataModule.SynchronizeAction  TTBXItem
TBXItem156Action)NonVisualDataModule.FullSynchronizeActionDisplayModenbdmImageAndText  TTBXSeparatorItemTBXSeparatorItem41  TTBXItem
TBXItem157Action!NonVisualDataModule.ConsoleAction  TTBXItem
TBXItem190ActionNonVisualDataModule.PuttyAction  TTBXSeparatorItemTBXSeparatorItem42  TTBXItem
TBXItem158Action-NonVisualDataModule.SynchronizeBrowsingAction   TTBXToolbarUpdatesToolbarLeft Top� CaptionUppdateringarDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXSubmenuItemTBXSubmenuItem1Action%NonVisualDataModule.ShowUpdatesActionDropdownCombo	 TTBXItem
TBXItem184Action)NonVisualDataModule.CheckForUpdatesAction  TTBXSeparatorItemTBXSeparatorItem46  TTBXItem
TBXItem180Action"NonVisualDataModule.HomepageAction  TTBXItem
TBXItem187Action&NonVisualDataModule.DownloadPageAction  TTBXItem
TBXItem181Action#NonVisualDataModule.ForumPageAction  TTBXItem
TBXItem182Action%NonVisualDataModule.HistoryPageAction  TTBXItem
TBXItem185Action$NonVisualDataModule.DonatePageAction  TTBXSeparatorItemTBXSeparatorItem45  TTBXItem
TBXItem183Action,NonVisualDataModule.UpdatesPreferencesAction    TTBXToolbarTransferToolbarLeft,Top� Caption   ÖverföringsinställningarDockPos,DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXLabelItemTransferSettingsLabelItemCaption   ÖverföringsinställningarMargin  TTBXDropDownItemTransferDropDown	EditWidth� Hint0   Välj förinställda överföringsinställningarDropDownList	 TTBXStringListTransferListMaxVisibleItemsMinWidth^  TTBXLabelItemTransferLabelMarginShowAccelChar  TTBXSeparatorItemTBXSeparatorItem52  TTBXItem
TBXItem189Action,NonVisualDataModule.PresetsPreferencesActionDisplayModenbdmImageAndText    TTBXToolbarCustomCommandsToolbarLeft+Top� CaptionEgna kommandonDockPos� DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrderVisible   �TPanelRemotePanelLeft�Top� Width�Height*Constraints.MinHeight� Constraints.MinWidth� TabOrder � 
TPathLabelRemotePathLabelLeft TopOWidth�HeightUnixPath	IndentVerticalAutoSizeVertical	HotTrack	OnGetStatusRemotePathLabelGetStatusOnPathClickRemotePathLabelPathClickAutoSizeTransparent
OnDblClickPathLabelDblClick  �	TSplitterRemotePanelSplitterLeft Top� Width�HeightCursorcrSizeNSHinti   Dra för att ändra storlek på katalogträd. Dubbelklicka för att gör höjden på katalogträden lika.AlignalTop  �TTBXStatusBarRemoteStatusBarTopWidth�SimplePanel	  �TUnixDirViewRemoteDirViewLeft Top� Width�Height|Constraints.MinHeightF
NortonLikenlOnOnUpdateStatusBarRemoteDirViewUpdateStatusBar	PathLabelRemotePathLabelAddParentDir	OnDDFileOperationExecuted(RemoteFileControlDDFileOperationExecutedOnHistoryGoDirViewHistoryGoOnPathChangeRemoteDirViewPathChange  �TUnixDriveViewRemoteDriveViewTopbWidth�Height-AlignalTopConstraints.MinHeightTabStop  TTBXDockRemoteTopDockLeft Top Width�HeightOColor	clBtnFaceFixAlign	 TTBXToolbarRemoteHistoryToolbarLeft TopCaption   FjärrhistorikDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXSubmenuItemRemoteBackButtonAction$NonVisualDataModule.RemoteBackActionDropdownCombo	  TTBXSubmenuItemRemoteForwardButtonAction'NonVisualDataModule.RemoteForwardActionDropdownCombo	   TTBXToolbarRemoteNavigationToolbarLeftFTopCaption   FjärrnavigeringDockPosDDockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem165Action)NonVisualDataModule.RemoteParentDirAction  TTBXItem
TBXItem166Action'NonVisualDataModule.RemoteRootDirAction  TTBXItem
TBXItem167Action'NonVisualDataModule.RemoteHomeDirAction  TTBXItem
TBXItem168Action'NonVisualDataModule.RemoteRefreshAction  TTBXSeparatorItemTBXSeparatorItem37  TTBXItem
TBXItem132Action)NonVisualDataModule.RemoteFindFilesActionDisplayModenbdmImageAndText  TTBXSeparatorItemTBXSeparatorItem44  TTBXItem
TBXItem170Action$NonVisualDataModule.RemoteTreeAction   TTBXToolbarRemotePathToolbarLeft Top Caption   Fjärrsökväg
DockableTodpTopdpBottom DockModedmCannotFloatDockPos ImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	Stretch	TabOrder OnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXComboBoxItemRemotePathComboBox	EditWidth� 	ShowImage	DropDownList	MaxVisibleItemsShowListImages	OnAdjustImageIndex"RemotePathComboBoxAdjustImageIndex
OnDrawItemRemotePathComboBoxDrawItemOnItemClickRemotePathComboBoxItemClickOnMeasureWidthRemotePathComboBoxMeasureWidthOnCancelRemotePathComboBoxCancel  TTBXItem
TBXItem169Action'NonVisualDataModule.RemoteOpenDirAction  TTBXItem
TBXItem229Action&NonVisualDataModule.RemoteFilterAction   TTBXToolbarRemoteFileToolbarLeftTop5Caption   FjärrfilerDockPosDockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem238Action$NonVisualDataModule.RemoteCopyActionDisplayModenbdmImageAndText  TTBXItem
TBXItem239Action$NonVisualDataModule.RemoteMoveAction  TTBXSeparatorItemTBXSeparatorItem55  TTBXItem
TBXItem242Action$NonVisualDataModule.RemoteEditActionDisplayModenbdmImageAndText  TTBXItem
TBXItem241Action&NonVisualDataModule.RemoteDeleteAction  TTBXItem
TBXItem240Action&NonVisualDataModule.RemoteRenameAction  TTBXItem
TBXItem243Action*NonVisualDataModule.RemotePropertiesActionDisplayModenbdmImageAndText  TTBXSeparatorItemTBXSeparatorItem56  TTBXItem
TBXItem244Action)NonVisualDataModule.RemoteCreateDirAction  TTBXItem
TBXItem246Action+NonVisualDataModule.RemoteAddEditLinkAction   TTBXToolbarRemoteSelectionToolbarLeft[Top5Caption   FjärrmarkeringDockPos[DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem138Action&NonVisualDataModule.RemoteSelectAction  TTBXItem
TBXItem139Action(NonVisualDataModule.RemoteUnselectAction  TTBXItem
TBXItem140Action)NonVisualDataModule.RemoteSelectAllAction    TTBXDockRemoteBottomDockLeft TopWidth�Height	Color	clBtnFaceFixAlign	PositiondpBottom   �TPanel
QueuePanelTopWidth=HeighttTabOrder �
TPathLabel
QueueLabelWidth=  �	TListView
QueueView3Width=HeightGTabStop  �TTBXDock	QueueDockWidth=   �TThemePageControlSessionsPageControlTop� Width=  TPanel
LocalPanelLeft Top� Width�Height*AlignalLeft
BevelOuterbvNoneColorclWindowConstraints.MinHeight� Constraints.MinWidth� ParentBackgroundTabOrder  
TPathLabelLocalPathLabelLeft TopOWidth�HeightIndentVerticalAutoSizeVertical	HotTrack	OnGetStatusLocalPathLabelGetStatusOnPathClickLocalPathLabelPathClickAutoSize	PopupMenu#NonVisualDataModule.LocalPanelPopupTransparent
OnDblClickPathLabelDblClick  	TSplitterLocalPanelSplitterLeft Top� Width�HeightCursorcrSizeNSHinti   Dra för att ändra storlek på katalogträd. Dubbelklicka för att gör höjden på katalogträden lika.AlignalTopAutoSnapColor	clBtnFaceMinSizeFParentColorResizeStylersUpdate  TTBXStatusBarLocalStatusBarLeft TopWidth�HeightPanels ParentShowHintSimplePanel	ShowHint	UseSystemFontOnClickLocalStatusBarClick  TDirViewLocalDirViewLeft Top� Width�Height|AlignalClientConstraints.MinHeightFDoubleBuffered	FullDrag	HideSelectionParentDoubleBuffered	PopupMenu%NonVisualDataModule.LocalDirViewPopupTabOrder	ViewStylevsReportOnColumnRightClickDirViewColumnRightClick	OnEditingDirViewEditingOnEnterLocalDirViewEnterDirColProperties.ExtVisible	PathLabelLocalPathLabelOnUpdateStatusBarLocalDirViewUpdateStatusBarOnGetSelectFilterRemoteDirViewGetSelectFilterHeaderImagesGlyphsModule.ArrowImagesAddParentDir	OnSelectItemDirViewSelectItemOnLoadedDirViewLoadedOnDDDragEnterLocalFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDDragOverLocalFileControlDDDragOverOnDDTargetHasDropHandler"LocalDirViewDDTargetHasDropHandlerOnDDFileOperationLocalFileControlDDFileOperationOnDDMenuPopupLocalFileControlDDMenuPopup
OnExecFileLocalDirViewExecFileOnMatchMaskDirViewMatchMaskOnGetOverlayDirViewGetOverlayConfirmDeleteWatchForChanges	OnFileIconForNameLocalDirViewFileIconForNameOnContextPopupLocalDirViewContextPopupOnHistoryChangeDirViewHistoryChangeOnHistoryGoDirViewHistoryGoOnPathChangeLocalDirViewPathChange  TTBXDockLocalTopDockLeft Top Width�HeightOColor	clBtnFaceFixAlign	 TTBXToolbarLocalHistoryToolbarLeft TopCaptionLokal historikDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXSubmenuItemLocalBackButtonAction#NonVisualDataModule.LocalBackActionDropdownCombo	  TTBXSubmenuItemLocalForwardButtonAction&NonVisualDataModule.LocalForwardActionDropdownCombo	   TTBXToolbarLocalNavigationToolbarLeftFTopCaptionLokal navigeringDockPosDDockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem159Action(NonVisualDataModule.LocalParentDirAction  TTBXItem
TBXItem160Action&NonVisualDataModule.LocalRootDirAction  TTBXItem
TBXItem161Action&NonVisualDataModule.LocalHomeDirAction  TTBXItem
TBXItem162Action&NonVisualDataModule.LocalRefreshAction  TTBXSeparatorItemTBXSeparatorItem43  TTBXItem
TBXItem164Action#NonVisualDataModule.LocalTreeAction   TTBXToolbarLocalPathToolbarLeft Top Caption   Lokal sökväg
DockableTodpTopdpBottom DockModedmCannotFloatDockPos ImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	Stretch	TabOrder OnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXComboBoxItemLocalPathComboBox	EditWidth� 	ShowImage	DropDownList	MaxVisibleItemsShowListImages	OnAdjustImageIndex!LocalPathComboBoxAdjustImageIndexOnItemClickLocalPathComboBoxItemClickOnCancelLocalPathComboBoxCancel  TTBXItem
TBXItem163Action&NonVisualDataModule.LocalOpenDirAction  TTBXItem
TBXItem228Action%NonVisualDataModule.LocalFilterAction   TTBXToolbarLocalFileToolbarLeft Top5CaptionLokala filerDockPos DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem231Action#NonVisualDataModule.LocalCopyActionDisplayModenbdmImageAndText  TTBXItem
TBXItem232Action#NonVisualDataModule.LocalMoveAction  TTBXSeparatorItemTBXSeparatorItem54  TTBXItem
TBXItem235Action#NonVisualDataModule.LocalEditActionDisplayModenbdmImageAndText  TTBXItem
TBXItem234Action%NonVisualDataModule.LocalDeleteAction  TTBXItem
TBXItem233Action%NonVisualDataModule.LocalRenameAction  TTBXItem
TBXItem236Action)NonVisualDataModule.LocalPropertiesActionDisplayModenbdmImageAndText  TTBXSeparatorItemTBXSeparatorItem35  TTBXItem
TBXItem237Action(NonVisualDataModule.LocalCreateDirAction  TTBXItem
TBXItem245Action*NonVisualDataModule.LocalAddEditLinkAction   TTBXToolbarLocalSelectionToolbarLeftITop5CaptionLokal markeringDockPosIDockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem137Action%NonVisualDataModule.LocalSelectAction  TTBXItem	TBXItem32Action'NonVisualDataModule.LocalUnselectAction  TTBXItem	TBXItem30Action(NonVisualDataModule.LocalSelectAllAction    
TDriveViewLocalDriveViewLeft TopbWidth�Height-WatchDirectory	DirViewLocalDirViewOnRefreshDrivesLocalDriveViewRefreshDrivesOnDDDragEnterLocalFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDDragOverLocalFileControlDDDragOverOnDDFileOperationLocalFileControlDDFileOperationOnDDMenuPopupLocalFileControlDDMenuPopupAlignalTopConstraints.MinHeightDoubleBuffered	HideSelectionIndentParentColorParentDoubleBufferedTabOrderTabStopOnEnterLocalDriveViewEnter  TTBXDockLocalBottomDockLeft TopWidth�Height	Color	clBtnFaceFixAlign	PositiondpBottom   TTBXDock
BottomDockLeft Top�Width=Height5FixAlign	PositiondpBottom TTBXToolbarToolbar2ToolbarLeft TopCaptionSnabbtangenterDockPos DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHintStretch	TabOrder Visible TTBXItem
TBXItem171Action'NonVisualDataModule.CurrentRenameActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem172Action%NonVisualDataModule.CurrentEditActionDisplayModenbdmImageAndTextStretch	  TTBXItemCurrentCopyToolbar2ItemAction$NonVisualDataModule.RemoteCopyActionDisplayModenbdmImageAndTextStretch	  TTBXItemCurrentMoveToolbar2ItemAction$NonVisualDataModule.RemoteMoveActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem175Action*NonVisualDataModule.CurrentCreateDirActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem176Action'NonVisualDataModule.CurrentDeleteActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem177Action+NonVisualDataModule.CurrentPropertiesActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem178Action*NonVisualDataModule.CloseApplicationActionDisplayModenbdmImageAndText
ImageIndex=Stretch	   TTBXToolbarCommandLineToolbarLeft Top CaptionCommandLineToolbarDockModedmCannotFloatStretch	TabOrderVisibleOnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXLabelItemCommandLinePromptLabelCaption
CommandX >Margin  TTBXComboBoxItemCommandLineComboOnBeginEditCommandLineComboBeginEditExtendedAccept	OnPopupCommandLineComboPopup    TTBXStatusBar	StatusBarLeft Top�Width=ImagesGlyphsModule.SessionImagesPanelsSizedStretchPriorityTag TextTruncationtwEndEllipsis 	AlignmenttaCenter
ImageIndexMaxSize#Size#Tag  	AlignmenttaCenterMaxSizeFViewPrioritybSizeFTag TextTruncationtwEndEllipsis 	AlignmenttaCenter
ImageIndex MaxSize#Size#Tag  	AlignmenttaCenterMaxSizePViewPrioritycSizePTag TextTruncationtwEndEllipsis  ParentShowHint	PopupMenu%NonVisualDataModule.CommanderBarPopupShowHint	UseSystemFontOnPanelDblClickStatusBarPanelDblClick  TPanelQueueSeparatorPanelLeft TopWidth=HeightAlignalBottom
BevelEdgesbeBottom 	BevelKindbkFlatTabOrder      TPF0�TScpExplorerFormScpExplorerFormLeft� Top� HelpType	htKeywordHelpKeywordui_explorerActiveControlRemoteDirViewCaptionScpExplorerFormClientHeight�ClientWidthxOldCreateOrder	PixelsPerInch`
TextHeight �	TSplitterQueueSplitterTopLWidthx  �TTBXDockTopDockWidthxHeight�  TTBXToolbarMenuToolbarLeft Top CaptionMenyCloseButtonImagesGlyphsModule.ExplorerImagesMenuBar	
ShrinkModetbsmWrapStretch	TabOrder  TTBXSubmenuItemTBXSubmenuItem5Caption&FilHelpKeywordui_explorer_menu#fileHintFiloperationer TTBXSubmenuItemTBXSubmenuItem26Caption&NyHelpKeyword
task_indexHintSkapa objekt|Skapa nytt objekt TTBXItem
TBXItem135Action!NonVisualDataModule.NewFileAction  TTBXItem
TBXItem136Action NonVisualDataModule.NewDirAction  TTBXItem
TBXItem209Action!NonVisualDataModule.NewLinkAction   TTBXSeparatorItemTBXSeparatorItem20  TTBXItem	TBXItem25Action%NonVisualDataModule.CurrentOpenAction  TTBXItem	TBXItem26Action$NonVisualDataModule.RemoteEditAction  TTBXSubmenuItemTBXSubmenuItem9Action0NonVisualDataModule.CurrentEditAlternativeAction  TTBXItemTBXItem4Action+NonVisualDataModule.RemoteAddEditLinkAction  TTBXSeparatorItemTBXSeparatorItem7  TTBXItem	TBXItem34Action&NonVisualDataModule.RemoteDeleteAction  TTBXItem	TBXItem35Action&NonVisualDataModule.RemoteRenameAction  TTBXItem	TBXItem41Action*NonVisualDataModule.RemotePropertiesAction  TTBXSeparatorItemTBXSeparatorItem8  TTBXItem	TBXItem30Action$NonVisualDataModule.RemoteCopyAction  TTBXItem	TBXItem32Action$NonVisualDataModule.RemoteMoveAction  TTBXItem	TBXItem31Action&NonVisualDataModule.RemoteCopyToAction  TTBXItem	TBXItem33Action&NonVisualDataModule.RemoteMoveToAction  TTBXItem	TBXItem36ActionNonVisualDataModule.PasteAction  TTBXSeparatorItemTBXSeparatorItem9  TTBXSubmenuItemCustomCommandsMenuAction(NonVisualDataModule.CustomCommandsAction  TTBXSubmenuItemTBXSubmenuItem6Caption&FilnamnHelpKeyword	filenamesHint$   Operationer med namn på valda filer TTBXItem	TBXItem38Action-NonVisualDataModule.FileListToClipboardAction  TTBXItem	TBXItem39Action1NonVisualDataModule.FullFileListToClipboardAction  TTBXItem	TBXItem40Action(NonVisualDataModule.UrlToClipboardAction   TTBXSeparatorItemTBXSeparatorItem1  TTBXItemTBXItem1Action&NonVisualDataModule.CloseSessionAction  TTBXItemTBXItem2Action*NonVisualDataModule.CloseApplicationAction   TTBXSubmenuItemTBXSubmenuItem7Caption
&KommandonHelpKeywordui_explorer_menu#commandsHintAndra kommandon TTBXItem	TBXItem43Action%NonVisualDataModule.SynchronizeAction  TTBXItem	TBXItem44Action)NonVisualDataModule.FullSynchronizeAction  TTBXItemTBXItem3Action)NonVisualDataModule.RemoteFindFilesAction  TTBXSubmenuItemQueueSubmenuItemCaption   &KöHelpKeywordui_queue#managing_the_queueHint   Kommandon för kölistaOnPopupQueueSubmenuItemPopup TTBXItemQueueEnableItem2Action%NonVisualDataModule.QueueEnableAction  TTBXItem	TBXItem46Action#NonVisualDataModule.QueueGoToAction  TTBXSeparatorItemTBXSeparatorItem10  TTBXItem	TBXItem47Action(NonVisualDataModule.QueueItemQueryAction  TTBXItem	TBXItem48Action(NonVisualDataModule.QueueItemErrorAction  TTBXItem	TBXItem49Action)NonVisualDataModule.QueueItemPromptAction  TTBXSeparatorItemTBXSeparatorItem11  TTBXItem	TBXItem50Action*NonVisualDataModule.QueueItemExecuteAction  TTBXItem
TBXItem196Action(NonVisualDataModule.QueueItemPauseAction  TTBXItem
TBXItem197Action)NonVisualDataModule.QueueItemResumeAction  TTBXItem	TBXItem51Action)NonVisualDataModule.QueueItemDeleteAction  TTBXComboBoxItemQueueSpeedComboBoxItemAction(NonVisualDataModule.QueueItemSpeedAction  TTBXSeparatorItemTBXSeparatorItem12  TTBXItem	TBXItem52Action%NonVisualDataModule.QueueItemUpAction  TTBXItem	TBXItem53Action'NonVisualDataModule.QueueItemDownAction  TTBXSeparatorItemTBXSeparatorItem48  TTBXSubmenuItemTBXSubmenuItem13Caption&AllaHelpKeywordui_queue#managing_the_queueHint&   Administrationskommandon för kömassa TTBXItem
TBXItem198Action'NonVisualDataModule.QueuePauseAllAction  TTBXItem
TBXItem199Action(NonVisualDataModule.QueueResumeAllAction  TTBXSeparatorItemTBXSeparatorItem35  TTBXItem
TBXItem143Action,NonVisualDataModule.QueueDeleteAllDoneAction    TTBXSeparatorItemTBXSeparatorItem13  TTBXItemTBXItem5Action+NonVisualDataModule.RemoteAddBookmarkAction  TTBXItemTBXItem6Action/NonVisualDataModule.RemotePathToClipboardAction  TTBXSeparatorItemTBXSeparatorItem2  TTBXItem	TBXItem54Action!NonVisualDataModule.ConsoleAction  TTBXItem	TBXItem55ActionNonVisualDataModule.PuttyAction  TTBXSeparatorItemTBXSeparatorItem14  TTBXItem	TBXItem56Action(NonVisualDataModule.FileSystemInfoAction  TTBXItem	TBXItem57Action%NonVisualDataModule.ClearCachesAction   TTBXSubmenuItemTBXSubmenuItem18Caption&MarkeraHelpKeywordui_explorer_menu#markHint   Kommandon för markera TTBXItem
TBXItem107Action#NonVisualDataModule.SelectOneAction  TTBXItem
TBXItem108Action NonVisualDataModule.SelectAction  TTBXItem
TBXItem109Action"NonVisualDataModule.UnselectAction  TTBXItem
TBXItem110Action#NonVisualDataModule.SelectAllAction  TTBXItem
TBXItem111Action)NonVisualDataModule.InvertSelectionAction  TTBXItem
TBXItem112Action(NonVisualDataModule.ClearSelectionAction  TTBXItem	TBXItem27Action*NonVisualDataModule.RestoreSelectionAction   TTBXSubmenuItemTBXSubmenuItem19CaptionSessionHelpKeywordui_explorer_menu#sessionHint   Kommandon för session TTBXItem
TBXItem113Action$NonVisualDataModule.NewSessionAction  TTBXItem	TBXItem90Action*NonVisualDataModule.DuplicateSessionAction  TTBXItem
TBXItem115Action&NonVisualDataModule.CloseSessionAction  TTBXItem
TBXItem114Action-NonVisualDataModule.SaveCurrentSessionAction2  TTBXSeparatorItemTBXSeparatorItem29  TTBXSubmenuItemTBXSubmenuItem21Action(NonVisualDataModule.OpenedSessionsAction  TTBXSubmenuItemTBXSubmenuItem231Action$NonVisualDataModule.WorkspacesAction  TTBXItem
TBXItem230Action'NonVisualDataModule.SaveWorkspaceAction  TTBXSeparatorItemTBXSeparatorItem53  TTBXSubmenuItemTBXSubmenuItem20Action(NonVisualDataModule.SavedSessionsAction2   TTBXSubmenuItemTBXSubmenuItem1Caption&VisaHelpKeywordui_explorer_menu#viewHint   Ändra layout för program TTBXSubmenuItemTBXSubmenuItem2Caption   &VerktygsfältHelpKeywordui_toolbarsHint   Visa/dölj verktygsfält TTBXItemTBXItem7Action-NonVisualDataModule.ExplorerAddressBandAction  TTBXItemTBXItem8Action-NonVisualDataModule.ExplorerToolbarBandAction  TTBXItemTBXItem9Action/NonVisualDataModule.ExplorerSelectionBandAction  TTBXItem	TBXItem10Action-NonVisualDataModule.ExplorerSessionBandAction  TTBXItem	TBXItem11Action1NonVisualDataModule.ExplorerPreferencesBandAction  TTBXItem	TBXItem12Action*NonVisualDataModule.ExplorerSortBandAction  TTBXItem	TBXItem82Action-NonVisualDataModule.ExplorerUpdatesBandAction  TTBXItem	TBXItem83Action.NonVisualDataModule.ExplorerTransferBandAction  TTBXItem	TBXItem28Action4NonVisualDataModule.ExplorerCustomCommandsBandAction  TTBXSeparatorItemTBXSeparatorItem19  TTBXItem	TBXItem92Action&NonVisualDataModule.LockToolbarsAction  TTBXItem
TBXItem140Action.NonVisualDataModule.SelectiveToolbarTextAction   TTBXItemSessionsTabsAction3Action&NonVisualDataModule.SessionsTabsAction  TTBXItem	TBXItem13Action#NonVisualDataModule.StatusBarAction  TTBXItem	TBXItem14Action!NonVisualDataModule.ViewLogAction  TTBXSubmenuItemTBXSubmenuItem14Caption   &KöHelpKeywordui_queueHint   Konfigurera kölista TTBXItem	TBXItem77Action#NonVisualDataModule.QueueShowAction	RadioItem	  TTBXItem	TBXItem78Action,NonVisualDataModule.QueueHideWhenEmptyAction	RadioItem	  TTBXItem	TBXItem79Action#NonVisualDataModule.QueueHideAction	RadioItem	  TTBXSeparatorItemTBXSeparatorItem21  TTBXItem	TBXItem80Action&NonVisualDataModule.QueueToolbarAction  TTBXSeparatorItemTBXSeparatorItem22  TTBXSubmenuItemTBXSubmenuItem8Action-NonVisualDataModule.QueueCycleOnceEmptyActionDropdownCombo	 TTBXItem
TBXItem222Action,NonVisualDataModule.QueueIdleOnceEmptyAction	RadioItem	  TTBXItem
TBXItem223Action2NonVisualDataModule.QueueDisconnectOnceEmptyAction	RadioItem	  TTBXItem
TBXItem224Action0NonVisualDataModule.QueueShutDownOnceEmptyAction	RadioItem	   TTBXItem	TBXItem81Action*NonVisualDataModule.QueuePreferencesAction   TTBXItem	TBXItem15Action$NonVisualDataModule.RemoteTreeAction  TTBXSeparatorItemTBXSeparatorItem3  TTBXItem	TBXItem16Action%NonVisualDataModule.CurrentIconAction  TTBXItem	TBXItem17Action*NonVisualDataModule.CurrentSmallIconAction  TTBXItem	TBXItem18Action%NonVisualDataModule.CurrentListAction  TTBXItem	TBXItem19Action'NonVisualDataModule.CurrentReportAction  TTBXSeparatorItemTBXSeparatorItem4  TTBXSubmenuItemTBXSubmenuItem15Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItem	TBXItem84Action'NonVisualDataModule.RemoteOpenDirAction  TTBXSeparatorItemTBXSeparatorItem25  TTBXItem	TBXItem85Action)NonVisualDataModule.RemoteParentDirAction  TTBXItem	TBXItem86Action'NonVisualDataModule.RemoteRootDirAction  TTBXItem	TBXItem87Action'NonVisualDataModule.RemoteHomeDirAction  TTBXSeparatorItemTBXSeparatorItem26  TTBXItem	TBXItem88Action$NonVisualDataModule.RemoteBackAction  TTBXItem	TBXItem89Action'NonVisualDataModule.RemoteForwardAction   TTBXItem	TBXItem20Action'NonVisualDataModule.RemoteRefreshAction  TTBXSubmenuItemTBXSubmenuItem16Caption&SorteraHelpKeywordui_file_panel#sorting_filesHint   Ändra filordning i panelen TTBXItem	TBXItem93Action-NonVisualDataModule.RemoteSortAscendingAction  TTBXSeparatorItemTBXSeparatorItem28  TTBXItem	TBXItem94Action*NonVisualDataModule.RemoteSortByNameAction
GroupIndex  TTBXItem	TBXItem95Action)NonVisualDataModule.RemoteSortByExtAction
GroupIndex  TTBXItem
TBXItem132Action*NonVisualDataModule.RemoteSortByTypeAction	RadioItem	  TTBXItem	TBXItem96Action-NonVisualDataModule.RemoteSortByChangedAction
GroupIndex  TTBXItem	TBXItem97Action*NonVisualDataModule.RemoteSortBySizeAction
GroupIndex  TTBXItem	TBXItem98Action,NonVisualDataModule.RemoteSortByRightsAction
GroupIndex  TTBXItem	TBXItem99Action+NonVisualDataModule.RemoteSortByOwnerAction
GroupIndex  TTBXItem
TBXItem100Action+NonVisualDataModule.RemoteSortByGroupAction
GroupIndex   TTBXSubmenuItemTBXSubmenuItem17CaptionVisa &kolumnerHelpKeywordui_file_panel#selecting_columnsHint$   Välj kolumner som ska visas i panel TTBXItem
TBXItem101Action2NonVisualDataModule.ShowHideRemoteNameColumnAction  TTBXItem
TBXItem102Action2NonVisualDataModule.ShowHideRemoteSizeColumnAction  TTBXItem
TBXItem131Action2NonVisualDataModule.ShowHideRemoteTypeColumnAction  TTBXItem
TBXItem103Action5NonVisualDataModule.ShowHideRemoteChangedColumnAction  TTBXItem
TBXItem104Action4NonVisualDataModule.ShowHideRemoteRightsColumnAction  TTBXItem
TBXItem105Action3NonVisualDataModule.ShowHideRemoteOwnerColumnAction  TTBXItem
TBXItem106Action3NonVisualDataModule.ShowHideRemoteGroupColumnAction  TTBXItem	TBXItem76Action8NonVisualDataModule.ShowHideRemoteLinkTargetColumnAction   TTBXItem
TBXItem138Action&NonVisualDataModule.RemoteFilterAction  TTBXSeparatorItemTBXSeparatorItem23  TTBXColorItemColorMenuItemAction#NonVisualDataModule.ColorMenuActionColorclNone  TTBXSeparatorItemTBXSeparatorItem5  TTBXItem	TBXItem21Action%NonVisualDataModule.PreferencesAction   TTBXSubmenuItemTBXSubmenuItem22Caption   &HjälpHelpKeywordui_explorer_menu#helpHint   Hjälp TTBXItem
TBXItem116Action)NonVisualDataModule.TableOfContentsAction  TTBXSeparatorItemTBXSeparatorItem30  TTBXItem
TBXItem117Action"NonVisualDataModule.HomepageAction  TTBXItem
TBXItem118Action#NonVisualDataModule.ForumPageAction  TTBXItem
TBXItem119Action%NonVisualDataModule.HistoryPageAction  TTBXSeparatorItemTBXSeparatorItem31  TTBXItem
TBXItem120Action)NonVisualDataModule.CheckForUpdatesAction  TTBXSeparatorItemTBXSeparatorItem32  TTBXItem
TBXItem121Action$NonVisualDataModule.DonatePageAction  TTBXSeparatorItemTBXSeparatorItem33  TTBXItem
TBXItem122ActionNonVisualDataModule.AboutAction    TTBXToolbarButtonsToolbarLeft Top4Caption	KommandonDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXSubmenuItem
BackButtonAction$NonVisualDataModule.RemoteBackActionDropdownCombo	  TTBXSubmenuItemForwardButtonAction'NonVisualDataModule.RemoteForwardActionDropdownCombo	  TTBXSeparatorItemTBXSeparatorItem6  TTBXItem	TBXItem23Action)NonVisualDataModule.RemoteParentDirAction  TTBXItem	TBXItem24Action'NonVisualDataModule.RemoteRootDirAction  TTBXItem	TBXItem29Action'NonVisualDataModule.RemoteHomeDirAction  TTBXItem	TBXItem37Action'NonVisualDataModule.RemoteRefreshAction  TTBXSeparatorItemTBXSeparatorItem24  TTBXItem
TBXItem139Action)NonVisualDataModule.RemoteFindFilesActionDisplayModenbdmImageAndText  TTBXSeparatorItemTBXSeparatorItem15  TTBXItem
TBXItem141Action$NonVisualDataModule.RemoteCopyActionDisplayModenbdmImageAndText  TTBXItem
TBXItem142Action$NonVisualDataModule.RemoteMoveAction  TTBXSeparatorItemTBXSeparatorItem27  TTBXItem	TBXItem42Action$NonVisualDataModule.RemoteEditActionDisplayModenbdmImageAndText  TTBXItem	TBXItem45Action%NonVisualDataModule.CurrentOpenAction  TTBXItem	TBXItem58Action&NonVisualDataModule.RemoteDeleteAction  TTBXItem	TBXItem59Action*NonVisualDataModule.RemotePropertiesActionDisplayModenbdmImageAndText  TTBXItem	TBXItem60Action&NonVisualDataModule.RemoteRenameAction  TTBXSeparatorItemTBXSeparatorItem16  TTBXItem	TBXItem61Action)NonVisualDataModule.RemoteCreateDirAction  TTBXItem	TBXItem62Action+NonVisualDataModule.RemoteAddEditLinkAction  TTBXItem	TBXItem63Action!NonVisualDataModule.ConsoleAction  TTBXItem	TBXItem91ActionNonVisualDataModule.PuttyAction  TTBXSeparatorItemTBXSeparatorItem17  TTBXItem	TBXItem64Action%NonVisualDataModule.SynchronizeAction  TTBXItem	TBXItem65Action)NonVisualDataModule.FullSynchronizeActionDisplayModenbdmImageAndText   TTBXToolbarSelectionToolbarLeft TopNCaption	MarkeringDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem	TBXItem66Action NonVisualDataModule.SelectAction  TTBXItem	TBXItem67Action"NonVisualDataModule.UnselectAction  TTBXSeparatorItemTBXSeparatorItem18  TTBXItem	TBXItem68Action#NonVisualDataModule.SelectAllAction  TTBXItem	TBXItem69Action)NonVisualDataModule.InvertSelectionAction  TTBXItem	TBXItem70Action(NonVisualDataModule.ClearSelectionAction  TTBXItem
TBXItem134Action*NonVisualDataModule.RestoreSelectionAction   TTBXToolbarSessionToolbarLeft TophCaptionSessionDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem123Action$NonVisualDataModule.NewSessionActionDisplayModenbdmImageAndText  TTBXItem
TBXItem137Action*NonVisualDataModule.DuplicateSessionAction  TTBXItem
TBXItem124Action&NonVisualDataModule.CloseSessionAction  TTBXItem
TBXItem125Action-NonVisualDataModule.SaveCurrentSessionAction2  TTBXSeparatorItemTBXSeparatorItem34  TTBXSubmenuItemTBXSubmenuItem23Action(NonVisualDataModule.SavedSessionsAction2DisplayModenbdmImageAndTextOptionstboDropdownArrow    TTBXToolbarPreferencesToolbarLeft Top� Caption   InställningarDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem126Action%NonVisualDataModule.PreferencesAction  TTBXSeparatorItemTBXSeparatorItem36  TTBXSubmenuItemTBXSubmenuItem3Action+NonVisualDataModule.CurrentCycleStyleActionDropdownCombo	 TTBXItem	TBXItem72Action%NonVisualDataModule.CurrentIconAction  TTBXItem	TBXItem73Action*NonVisualDataModule.CurrentSmallIconAction  TTBXItem	TBXItem74Action%NonVisualDataModule.CurrentListAction  TTBXItem	TBXItem75Action'NonVisualDataModule.CurrentReportAction   TTBXItem
TBXItem127Action!NonVisualDataModule.ViewLogAction  TTBXSubmenuItemTBXSubmenuItem24Action)NonVisualDataModule.QueueToggleShowActionDisplayModenbdmImageAndTextDropdownCombo	 TTBXItem
TBXItem128Action#NonVisualDataModule.QueueShowAction	RadioItem	  TTBXItem
TBXItem129Action,NonVisualDataModule.QueueHideWhenEmptyAction	RadioItem	  TTBXItem
TBXItem130Action#NonVisualDataModule.QueueHideAction	RadioItem	   TTBXItem	TBXItem71Action$NonVisualDataModule.RemoteTreeAction   TTBXToolbarSortToolbarLeft Top� CaptionSorteraDockPos DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXItem
TBXItem145Action.NonVisualDataModule.CurrentSortAscendingAction  TTBXSeparatorItemTBXSeparatorItem40  TTBXItem
TBXItem146Action+NonVisualDataModule.CurrentSortByNameAction  TTBXItem
TBXItem147Action*NonVisualDataModule.CurrentSortByExtAction  TTBXItem
TBXItem133Action*NonVisualDataModule.RemoteSortByTypeAction	RadioItem	  TTBXItem
TBXItem149Action.NonVisualDataModule.CurrentSortByChangedAction  TTBXItem
TBXItem150Action+NonVisualDataModule.CurrentSortBySizeAction  TTBXItem
TBXItem151Action-NonVisualDataModule.CurrentSortByRightsAction  TTBXItem
TBXItem152Action,NonVisualDataModule.CurrentSortByOwnerAction  TTBXItem
TBXItem153Action,NonVisualDataModule.CurrentSortByGroupAction   TTBXToolbarAddressToolbarLeft TopCaptionAdress
DockableTodpTopdpBottom DockModedmCannotFloatDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHint	PopupMenu&NonVisualDataModule.RemoteAddressPopup	ResizableShowHint	Stretch	TabOrderOnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXLabelItemTBXLabelItem1CaptionAdressMargin  TTBXComboBoxItemUnixPathComboBox	EditWidth� OnAcceptTextUnixPathComboBoxAcceptTextOnBeginEditUnixPathComboBoxBeginEdit	ShowImage	MaxVisibleItemsShowListImages	OnAdjustImageIndex"RemotePathComboBoxAdjustImageIndex
OnDrawItemRemotePathComboBoxDrawItemOnItemClickRemotePathComboBoxItemClickOnMeasureWidthRemotePathComboBoxMeasureWidthOnCancelRemotePathComboBoxCancel  TTBXItem	TBXItem22Action'NonVisualDataModule.RemoteOpenDirAction  TTBXItem
TBXItem229Action&NonVisualDataModule.RemoteFilterAction   TTBXToolbarUpdatesToolbarLeft Top� CaptionUppdateringarDockPos�DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXSubmenuItemTBXSubmenuItem4Action%NonVisualDataModule.ShowUpdatesActionDropdownCombo	 TTBXItem
TBXItem184Action)NonVisualDataModule.CheckForUpdatesAction  TTBXSeparatorItemTBXSeparatorItem46  TTBXItem
TBXItem180Action"NonVisualDataModule.HomepageAction  TTBXItem
TBXItem187Action&NonVisualDataModule.DownloadPageAction  TTBXItem
TBXItem181Action#NonVisualDataModule.ForumPageAction  TTBXItem
TBXItem182Action%NonVisualDataModule.HistoryPageAction  TTBXItem
TBXItem185Action$NonVisualDataModule.DonatePageAction  TTBXSeparatorItemTBXSeparatorItem45  TTBXItem
TBXItem183Action,NonVisualDataModule.UpdatesPreferencesAction    TTBXToolbarTransferToolbarLeft,Top� Caption   ÖverföringsinställningarDockPos,DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder TTBXLabelItemTransferSettingsLabelItemCaption   ÖverföringsinställningarMargin  TTBXDropDownItemTransferDropDown	EditWidth� Hint0   Välj förinställda överföringsinställningarDropDownList	 TTBXStringListTransferListMaxVisibleItemsMinWidth^  TTBXLabelItemTransferLabelMarginShowAccelChar  TTBXSeparatorItemTBXSeparatorItem52  TTBXItem
TBXItem189Action,NonVisualDataModule.PresetsPreferencesActionDisplayModenbdmImageAndText    TTBXToolbarCustomCommandsToolbarLeft+Top� CaptionEgna kommandonDockPos� DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder	Visible   �TPanelRemotePanelLeft	Top� WidthfHeightfConstraints.MinHeightdConstraints.MinWidth�  �	TSplitterRemotePanelSplitterHeightGHintW   Dra för att ändra storlek på katalogträd. Dubbelklicka för att dölja katalogträd  �TTBXStatusBarRemoteStatusBarTopPWidthfHeightImagesGlyphsModule.SessionImagesPanelsSizedStretchPriorityTag TextTruncationtwEndEllipsis 	AlignmenttaCenter
ImageIndexMaxSize#Size#Tag  	AlignmenttaCenterMaxSizeFViewPrioritybSizeFTag TextTruncationtwEndEllipsis 	AlignmenttaCenter
ImageIndex MaxSize#Size#Tag  	AlignmenttaCenterMaxSizePViewPrioritycSizePTag TextTruncationtwEndEllipsis  OnPanelDblClickStatusBarPanelDblClick  �TUnixDirViewRemoteDirViewWidth�HeightGOnUpdateStatusBarRemoteDirViewUpdateStatusBarOnPathChangeRemoteDirViewPathChange  �TUnixDriveViewRemoteDriveViewHeightGConstraints.MinWidth(  TTBXDock
BottomDockLeft TopGWidthfHeight	Color	clBtnFaceFixAlign	PositiondpBottom   �TPanel
QueuePanelTopOWidthx �
TPathLabel
QueueLabelWidthx  �	TListView
QueueView3Widthx  �TTBXDock	QueueDockWidthx   �TThemePageControlSessionsPageControlTop� Widthx  TTBXDockLeftDockLeft Top� Width	HeightfPositiondpLeft  TTBXDock	RightDockLeftoTop� Width	HeightfPositiondpRight    TPF0TSelectMaskDialogSelectMaskDialogLeftqTopHelpType	htKeywordHelpKeyword	ui_selectBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSelectXClientHeight� ClientWidthiColor	clBtnFace
ParentFont	OldCreateOrder	Position
poDesignedOnCloseQueryFormCloseQueryOnShowFormShow
DesignSizei�  PixelsPerInch`
TextHeight 	TGroupBox	MaskGroupLeftTopWidthYHeight^AnchorsakLeftakTopakRightakBottom TabOrder 
DesignSizeY^  TLabelLabel3LeftTopWidth/HeightCaption	Fil&mask:FocusControlMaskEdit  	TCheckBoxApplyToDirectoriesCheckLeftTop?Width� HeightCaption   Tillämpa på &katalogerTabOrder  THistoryComboBoxMaskEditLeftTop$Width9HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder Text*.*OnExitMaskEditExit  TStaticTextHintTextLeft� Top@WidthiHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	Mask&tipsTabOrderTabStop	   TButtonOKBtnLeftmTopmWidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft� TopmWidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeftTopmWidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TButtonClearButtonLeftTopmWidthKHeightAnchorsakRightakBottom Caption&RensaModalResultTabOrderOnClickClearButtonClick      TPF0TSiteAdvancedDialogSiteAdvancedDialogLeft_Top� HelpType	htKeywordHelpKeywordui_site_advancedBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption"   Avancerade webbplatsinställningarClientHeight�ClientWidth1Color	clBtnFace
ParentFont	OldCreateOrder	PositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize1� PixelsPerInch`
TextHeight TPanel	MainPanelLeft Top Width1Height�AlignalTopAnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneTabOrder  TPageControlPageControlTagLeft� Top Width�Height�HelpType	htKeyword
ActivePageEnvironmentSheetAlignalClient	MultiLine	Style	tsButtonsTabOrderTabStopOnChangePageControlChange 	TTabSheetEnvironmentSheetTagHelpType	htKeywordHelpKeywordui_login_environmentCaption   Miljö
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxEnvironmentGroupLeft TopWidth�Height`AnchorsakLeftakTopakRight Caption   ServermiljöTabOrder 
DesignSize�`  TLabelEOLTypeLabelLeftTopWidth� HeightCaption1   Slut på rad &tecken (om det inte ges av server):FocusControlEOLTypeCombo  TLabelUtfLabelLeftTop,Width� HeightCaption   &UTF-8 kodning på filnamn:FocusControlUtfCombo  TLabelTimeDifferenceLabelLeftTopDWidthQHeightCaptionOffset tidszon:FocusControlTimeDifferenceEdit  TLabelTimeDifferenceHoursLabelLeft� TopDWidthHeightAnchorsakTopakRight CaptiontimmarFocusControlTimeDifferenceEdit  TLabelTimeDifferenceMinutesLabelLeftPTopBWidth%HeightAnchorsakTopakRight CaptionminuterFocusControlTimeDifferenceMinutesEdit  	TComboBoxEOLTypeComboLeft@TopWidth=HeightStylecsDropDownListAnchorsakTopakRight TabOrder Items.StringsLFCR/LF   	TComboBoxUtfComboLeft@Top'Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrder  TUpDownEditTimeDifferenceEditLeft� Top?WidthEHeight	AlignmenttaRightJustifyMaxValue       �@MinValue       ��Value       ��AnchorsakTopakRight TabOrderOnChange
DataChange  TUpDownEditTimeDifferenceMinutesEditLeftTop?WidthEHeight	AlignmenttaRightJustify	Increment       �@MaxValue       �@MinValue       ��Value       ��AnchorsakTopakRight TabOrderOnChange
DataChange   	TGroupBoxDSTModeGroupLeft TopnWidth�Height]AnchorsakLeftakTopakRight Caption	SommartidTabOrder
DesignSize�]  TRadioButtonDSTModeUnixCheckLeftTopWidthqHeightAnchorsakLeftakTopakRight Caption7   Justera fjärrtidsstämpel med lokal ko&nvention (Unix)TabOrder OnClick
DataChange  TRadioButtonDSTModeWinCheckLeftTop*WidthqHeightAnchorsakLeftakTopakRight Caption-   Justera fjärrtidsstämpel med &DST (Windows)TabOrderOnClick
DataChange  TRadioButtonDSTModeKeepCheckLeftTopAWidthqHeightAnchorsakLeftakTopakRight Caption    Bevara fjärrtidsstämpel (Unix)TabOrderOnClick
DataChange    	TTabSheetDirectoriesSheetTagHelpType	htKeywordHelpKeywordui_login_directoriesCaption	Kataloger
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxDirectoriesGroupLeft TopWidth�Height� AnchorsakLeftakTopakRight Caption	KatalogerTabOrder 
DesignSize��   TLabelLocalDirectoryLabelLeftTopoWidthJHeightCaption&Lokal katalogFocusControlLocalDirectoryEdit  TLabelRemoteDirectoryLabelLeftTopBWidthWHeightCaption   F&järrkatalogFocusControlRemoteDirectoryEdit  TLabelLocalDirectoryDescLabelLeftTop� Width� HeightCaptionB   Lokal katalog används inte i det utforskar-liknande gränssnittet  TDirectoryEditLocalDirectoryEditLeftTop� WidthsHeightAcceptFiles	
DialogText    Välj lokal katalog vid uppstartClickKey@AnchorsakLeftakTopakRight TabOrderTextLocalDirectoryEditOnChange
DataChange  TEditRemoteDirectoryEditLeftTopSWidthsHeightAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRemoteDirectoryEditOnChange
DataChange  	TCheckBoxUpdateDirectoriesCheckLeftTop*WidthqHeightAnchorsakLeftakTopakRight Caption"   Ko&m ihåg senast använda katalogTabOrder  	TCheckBoxSynchronizeBrowsingCheckLeftTopWidthqHeightAnchorsakLeftakTopakRight Caption   Syn&kronisera bläddringTabOrder    	TGroupBoxDirectoryOptionsGroupLeft Top� Width�Height]AnchorsakLeftakTopakRight Caption   Alternativ vid kalalogläsningTabOrder
DesignSize�]  	TCheckBoxCacheDirectoriesCheckLeftTopWidthqHeightAnchorsakLeftakTopakRight Caption   Cacha &besökta fjärrkatalogerTabOrder OnClick
DataChange  	TCheckBoxCacheDirectoryChangesCheckLeftTop*Width� HeightAnchorsakLeftakTopakRight Caption   Cacha katalogf&örändringarTabOrderOnClick
DataChange  	TCheckBoxResolveSymlinksCheckLeftTopAWidthqHeightAnchorsakLeftakTopakRight Caption   Slå upp symboliska lä&nkarTabOrder  	TCheckBoxPreserveDirectoryChangesCheckLeft� Top*Width� HeightAnchorsakTopakRight Caption&Permanent cacheTabOrder    	TTabSheetRecycleBinSheetTagHelpType	htKeywordHelpKeywordui_login_recycle_binCaptionPapperskorg
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxRecycleBinGroupLeft TopWidth�HeightrAnchorsakLeftakTopakRight CaptionPapperskorgTabOrder 
DesignSize�r  TLabelRecycleBinPathLabelLeftTop@Width_HeightCaption   Papp&erskorg på servernFocusControlRecycleBinPathEdit  	TCheckBoxDeleteToRecycleBinCheckLeftTopWidthrHeightAnchorsakLeftakTopakRight Caption6   Flytta borttagna filer på servern till &papperskorgenTabOrder OnClick
DataChange  	TCheckBoxOverwrittenToRecycleBinCheckLeftTop*WidthrHeightAnchorsakLeftakTopakRight CaptionG   Flytta &överskrivna filer på servern till papperskorgen (endast SFTP)TabOrderOnClick
DataChange  TEditRecycleBinPathEditLeftTopQWidthrHeightAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRecycleBinPathEditOnChange
DataChange    	TTabSheet	SftpSheetTagHelpType	htKeywordHelpKeywordui_login_sftpCaptionSFTP
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxSFTPBugsGroupBoxLeft ToplWidth�HeightFAnchorsakLeftakTopakRight Caption    Upptäckta buggar i SFTP servrarTabOrder
DesignSize�F  TLabelLabel10LeftTopWidth� HeightCaption;   &Omvänd ordning på symboliska länkar i kommandoargument:FocusControlSFTPBugSymlinkCombo  TLabelLabel36LeftTop,Width� HeightCaption3   Feltolkning av filtidsstä&mplar tidigare än 1970:FocusControlSFTPBugSignedTSCombo  	TComboBoxSFTPBugSymlinkComboLeft@TopWidth=HeightStylecsDropDownListAnchorsakTopakRight TabOrder   	TComboBoxSFTPBugSignedTSComboLeft@Top'Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrder   	TGroupBoxSFTPProtocolGroupLeft TopWidth�Height`AnchorsakLeftakTopakRight Caption   Alternativ för protokollTabOrder 
DesignSize�`  TLabelLabel34LeftTop,Width� HeightCaption"   Före&drar SFTP protokoll version:FocusControlSFTPMaxVersionCombo  TLabelLabel23LeftTopWidth>HeightCaptionSFTP ser&verFocusControlSftpServerEdit  	TComboBoxSFTPMaxVersionComboLeft@Top'Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderItems.Strings012345   	TComboBoxSftpServerEditLeft� TopWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength� TabOrder TextSftpServerEditItems.StringsStandard/bin/sftp-serversudo su -c /bin/sftp-server   	TCheckBoxAllowScpFallbackCheckLeftTopDWidthqHeightAnchorsakLeftakTopakRight Caption   Tillåt SCP &fallbackTabOrderOnClick
DataChange    	TTabSheetScpSheetTagHelpType	htKeywordHelpKeywordui_login_scpCaption
SCP/ShellX
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxOtherShellOptionsGroupLeft Top� Width�HeightEAnchorsakLeftakTopakRight Caption   Övriga alternativTabOrder
DesignSize�E  	TCheckBoxLookupUserGroupsCheckLeftTopWidth� HeightAllowGrayed	Caption   Slå upp &användargrupperTabOrder OnClick
DataChange  	TCheckBoxClearAliasesCheckLeftTop*Width� HeightCaptionRensa a&liasTabOrderOnClick
DataChange  	TCheckBoxUnsetNationalVarsCheckLeft� TopWidth� HeightAnchorsakLeftakTopakRight CaptionRensa &nationella variablerTabOrderOnClick
DataChange  	TCheckBoxScp1CompatibilityCheckLeft� Top*Width� HeightAnchorsakLeftakTopakRight Caption%   Använd scp&2 med scp1 kompatibilitetTabOrderOnClick
DataChange   	TGroupBox
ShellGroupLeft TopWidth�HeightFAnchorsakLeftakTopakRight CaptionSkalTabOrder 
DesignSize�F  TLabelLabel19LeftTopWidthHeightCaptionS&kal:FocusControl	ShellEdit  TLabelLabel20LeftTop,WidthhHeightCaption&Returnera kodvariabel:FocusControlReturnVarEdit  	TComboBox	ShellEditLeft� TopWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength2TabOrder Text	ShellEditItems.StringsStandard	/bin/bash/bin/ksh	sudo su -   	TComboBoxReturnVarEditLeft� Top'Width� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength2TabOrderTextReturnVarEditItems.StringsDetektera automatiskt?status    	TGroupBoxScpLsOptionsGroupLeft TopTWidth�HeightEAnchorsakLeftakTopakRight CaptionListning av katalogerTabOrder
DesignSize�E  TLabelLabel9LeftTopWidthRHeightCaption   &Kommando för listning:FocusControlListingCommandEdit  	TCheckBoxIgnoreLsWarningsCheckLeftTop*Width� HeightCaptionIgnorera LS &varningarTabOrderOnClick
DataChange  	TCheckBoxSCPLsFullTimeAutoCheckLeft� Top*Width� HeightAnchorsakLeftakTopakRight Caption#   Försök att få &full tidsstämpelTabOrderOnClick
DataChange  	TComboBoxListingCommandEditLeft� TopWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength2TabOrder TextListingCommandEditItems.Stringsls -lals -gla     	TTabSheetFtpSheetTagHelpType	htKeywordHelpKeywordui_login_ftpCaptionFTP
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxFtpGroupLeft TopWidth�Height� AnchorsakLeftakTopakRight Caption   Alternativ för protokollTabOrder 
DesignSize��   TLabelLabel25LeftTop*WidthgHeightCaption&Kommandon efter inloggning:FocusControlPostLoginCommandsMemo  TLabelFtpListAllLabelLeftTop� Width� HeightCaption%   &Support för listning av dolda filerFocusControlFtpListAllCombo  TLabelLabel24LeftTop|Width� HeightCaption,   Använd &MLSD kommandon för kataloglistningFocusControlFtpUseMlsdCombo  TLabelFtpForcePasvIpLabelLeftTop� Width� HeightCaption+   &Tvinga ip-adress för passiva anslutningarFocusControlFtpForcePasvIpCombo  TLabelFtpAccountLabelLeftTopWidth+HeightCaptionK&onto:FocusControlFtpAccountEdit  TMemoPostLoginCommandsMemoLeftTop;WidthqHeight5AnchorsakLeftakTopakRight 
ScrollBars
ssVerticalTabOrder  	TComboBoxFtpListAllComboLeft@Top� Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxFtpForcePasvIpComboLeft@Top� Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxFtpUseMlsdComboLeft@TopwWidth=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  TEditFtpAccountEditLeft� TopWidth� HeightAnchorsakLeftakTopakRight 	MaxLengthdTabOrder TextFtpAccountEditOnChange
DataChange    	TTabSheet	ConnSheetTagHelpType	htKeywordHelpKeywordui_login_connectionCaption
Anslutning
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxFtpPingGroupLeft Top� Width�HeightuAnchorsakLeftakTopakRight Caption
KeepalivesTabOrder
DesignSize�u  TLabelFtpPingIntervalLabelLeftTopZWidth� HeightCaptionSekunder &mellan keepalivesFocusControlFtpPingIntervalSecEdit  TUpDownEditFtpPingIntervalSecEditLeft� TopUWidthIHeight	AlignmenttaRightJustifyMaxValue       �
@MinValue       ��?Value       ��?	MaxLengthTabOrderOnChange
DataChange  TRadioButtonFtpPingOffButtonLeftTopWidthmHeightAnchorsakLeftakTopakRight Caption&AvTabOrder OnClick
DataChange  TRadioButtonFtpPingNullPacketButtonLeftTop*WidthmHeightAnchorsakLeftakTopakRight CaptionSkicka SSH-&null-paketEnabledTabOrderOnClick
DataChange  TRadioButtonFtpPingDummyCommandButtonLeftTopAWidthmHeightAnchorsakLeftakTopakRight Caption#   Kör kommandon för &dummy-protkollTabOrderOnClick
DataChange   	TGroupBoxTimeoutGroupLeft TopPWidth�Height.AnchorsakLeftakTopakRight Caption	TimeouterTabOrder
DesignSize�.  TLabelLabel11LeftTopWidthzHeightCaption   Timeout för se&rversvar:FocusControlTimeoutEdit  TLabelLabel12LeftNTopWidth'HeightAnchorsakTopakRight CaptionsekunderFocusControlTimeoutEdit  TUpDownEditTimeoutEditLeft TopWidthIHeight	AlignmenttaRightJustify	Increment       �@MaxValue      ��@MinValue       �@Value       �@AnchorsakTopakRight 	MaxLengthTabOrder OnChange
DataChange   	TGroupBox	PingGroupLeft Top� Width�HeightuAnchorsakLeftakTopakRight Caption
KeepalivesTabOrder
DesignSize�u  TLabelPingIntervalLabelLeftTopZWidth� HeightCaptionSekunder &mellan keepalivesFocusControlPingIntervalSecEdit  TUpDownEditPingIntervalSecEditLeft TopUWidthIHeight	AlignmenttaRightJustifyMaxValue       �
@MinValue       ��?Value       ��?AnchorsakTopakRight 	MaxLengthTabOrderOnChange
DataChange  TRadioButtonPingOffButtonLeftTopWidthmHeightAnchorsakLeftakTopakRight CaptionA&vTabOrder OnClick
DataChange  TRadioButtonPingNullPacketButtonLeftTop*WidthmHeightAnchorsakLeftakTopakRight CaptionSkicka SSH-&null-paketTabOrderOnClick
DataChange  TRadioButtonPingDummyCommandButtonLeftTopAWidthmHeightAnchorsakLeftakTopakRight Caption%   Kör kommandon för &dummy-protokoll:TabOrderOnClick
DataChange   	TGroupBoxIPvGroupLeft Top� Width�Height.AnchorsakLeftakTopakRight Caption   Version för internetprotokollTabOrder TRadioButtonIPAutoButtonLeftTopWidtheHeightCaptionA&utomatiskTabOrder OnClick
DataChange  TRadioButton
IPv4ButtonLeft|TopWidtheHeightCaptionIPv&4TabOrderOnClick
DataChange  TRadioButton
IPv6ButtonLeft� TopWidtheHeightCaptionIPv&6TabOrderOnClick
DataChange   	TGroupBoxConnectionGroupLeft TopWidth�HeightEAnchorsakLeftakTopakRight Caption
AnslutningTabOrder 
DesignSize�E  	TCheckBoxFtpPasvModeCheckLeftTopWidthqHeightAnchorsakLeftakTopakRight Caption   &Passivt lägeTabOrder OnClick
DataChange  	TCheckBoxBufferSizeCheckLeftTop*WidthqHeightAnchorsakLeftakTopakRight Caption(   Optimera storlek på anslutnings&buffertTabOrderOnClick
DataChange    	TTabSheet
ProxySheetTagHelpType	htKeywordHelpKeywordui_login_proxyCaptionProxy
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxProxyTypeGroupLeft TopWidth�Height� AnchorsakLeftakTopakRight CaptionProxyTabOrder 
DesignSize��   TLabelProxyMethodLabelLeftTopWidth9HeightCaption&Typ av proxy:FocusControlSshProxyMethodCombo  TLabelProxyHostLabelLeftTop)WidthUHeightCaption   Pro&xyns värdnamn:FocusControlProxyHostEdit  TLabelProxyPortLabelLeftTop)Width?HeightAnchorsakTopakRight CaptionPo&rtnummer:FocusControlProxyPortEdit  TLabelProxyUsernameLabelLeftTopUWidth7HeightCaption   &Användarnamn:FocusControlProxyUsernameEdit  TLabelProxyPasswordLabelLeft� TopUWidth2HeightCaption   &Lösenord:FocusControlProxyPasswordEdit  	TComboBoxSshProxyMethodComboLeft� TopWidthnHeightStylecsDropDownListTabOrder OnChange
DataChangeItems.StringsIngenSOCKS4SOCKS5HTTPTelnetLokal   TUpDownEditProxyPortEditLeftTop:WidthbHeight	AlignmenttaRightJustifyMaxValue      ��@MinValue       ��?Value       ��?AnchorsakTopakRight TabOrderOnChange
DataChange  TEditProxyHostEditLeftTop:Width
HeightAnchorsakLeftakTopakRight 	MaxLength2TabOrderTextProxyHostEditOnChange
DataChange  TEditProxyUsernameEditLeftTopfWidth� Height	MaxLength2TabOrderTextProxyUsernameEditOnChange
DataChange  TPasswordEditProxyPasswordEditLeft� TopfWidth� HeightAnchorsakLeftakTopakRight 	MaxLength2TabOrderTextProxyPasswordEditOnChange
DataChange  	TComboBoxFtpProxyMethodComboLeft� TopWidth� HeightStylecsDropDownListAnchorsakLeftakTopakRight DropDownCountTabOrderOnChange
DataChangeItems.StringsIngenSOCKS4SOCKS5HTTP
SITE %host!USER %proxyuser, USER %user@%host
OPEN %hostUSER %proxyuser, USER %userUSER %user@%hostUSER %proxyuser@%hostUSER %user@%host %proxyuserUSER %user@%proxyuser@%host   	TComboBoxWebDavProxyMethodComboLeft� TopWidthnHeightStylecsDropDownListTabOrderOnChange
DataChangeItems.StringsIngenSOCKS4SOCKS5HTTP    	TGroupBoxProxySettingsGroupLeft Top� Width�Height� AnchorsakLeftakTopakRight Caption   Inställningar proxyTabOrder
DesignSize��   TLabelProxyTelnetCommandLabelLeftTopWidthRHeightCaptionTelnetko&mmando:FocusControlProxyTelnetCommandEdit  TLabelLabel17LeftTopcWidth� HeightCaption-   Låt &DNS-namnuppslagningar göras av proxyn:  TLabelProxyLocalCommandLabelLeftTopWidthkHeightCaptionLokalt proxyko&mmando:FocusControlProxyLocalCommandEdit  TEditProxyTelnetCommandEditLeftTop#WidthrHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder TextProxyTelnetCommandEditOnChange
DataChange  	TCheckBoxProxyLocalhostCheckLeftTopMWidthrHeightAnchorsakLeftakTopakRight Caption(   Låt lokala a&nslutningar gå via proxynTabOrder  	TComboBoxProxyDNSComboLeft� Top^Width� HeightStylecsDropDownListAnchorsakLeftakTopakRight TabOrderItems.Strings
AutomatiskNejJa   TEditProxyLocalCommandEditLeftTop#WidthHeightAnchorsakLeftakTopakRight TabOrderTextProxyLocalCommandEditOnChange
DataChange  TButtonProxyLocalCommandBrowseButtonLeft,Top!WidthRHeightAnchorsakTopakRight Caption   &Bläddra...TabOrderOnClick"ProxyLocalCommandBrowseButtonClick  TStaticTextProxyTelnetCommandHintTextLeft/Top:WidthOHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption   mönsterTabOrderTabStop	  TStaticTextProxyLocalCommandHintTextLeft� Top:WidthOHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption   mönsterTabOrderTabStop	    	TTabSheetTunnelSheetTagHelpType	htKeywordHelpKeywordui_login_tunnelCaptionTunnel
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxTunnelSessionGroupLeft Top Width�HeightvAnchorsakLeftakTopakRight Caption    Värd för att sätta upp tunnelTabOrder
DesignSize�v  TLabelLabel6LeftTopWidth7HeightCaption   &Värdnamn:FocusControlTunnelHostNameEdit  TLabelLabel14LeftTopWidth?HeightAnchorsakTopakRight CaptionPo&rtnummer:FocusControlTunnelPortNumberEdit  TLabelLabel15LeftTopDWidth7HeightCaption   &Användarnamn:FocusControlTunnelUserNameEdit  TLabelLabel16Left� TopDWidth2HeightCaption   &Lösenord:FocusControlTunnelPasswordEdit  TEditTunnelHostNameEditLeftTop#Width
HeightAnchorsakLeftakTopakRight 	MaxLengthdTabOrder TextTunnelHostNameEditOnChange
DataChange  TEditTunnelUserNameEditLeftTopUWidth� Height	MaxLength2TabOrderTextTunnelUserNameEditOnChange
DataChange  TPasswordEditTunnelPasswordEditLeft� TopUWidth� HeightAnchorsakLeftakTopakRight 	MaxLength2TabOrderTextTunnelPasswordEditOnChange
DataChange  TUpDownEditTunnelPortNumberEditLeftTop#WidthbHeight	AlignmenttaRightJustifyMaxValue      ��@MinValue       ��?Value       ��?AnchorsakTopakRight TabOrderOnChange
DataChange   	TCheckBoxTunnelCheckLeftTopWidth~HeightAnchorsakLeftakTopakRight CaptionAnslut med SSH-tunnelTabOrder OnClick
DataChange  	TGroupBoxTunnelOptionsGroupLeft Top� Width�Height/AnchorsakLeftakTopakRight Caption   Alternativ för tunnelTabOrder
DesignSize�/  TLabelLabel21LeftTopWidthTHeightCaption&Lokal tunnelport:FocusControlTunnelLocalPortNumberEdit  	TComboBoxTunnelLocalPortNumberEditLeftTopWidthbHeightAutoCompleteAnchorsakTopakRight 	MaxLength2TabOrder TextTunnelLocalPortNumberEditOnChange
DataChangeItems.Strings   Välj automatiskt    	TGroupBoxTunnelAuthenticationParamsGroupLeft Top� Width�HeightDAnchorsakLeftakTopakRight CaptionTunnelautentiseringsparametrarTabOrder
DesignSize�D  TLabelLabel18LeftTopWidthKHeightCaptionPrivat nyc&kelfilFocusControlTunnelPrivateKeyEdit  TFilenameEditTunnelPrivateKeyEditLeftTop#WidthrHeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPrivateKeyEditAfterDialogFilter8PuTTY privata nycklar (*.ppk)|*.ppk|Alla filer (*.*)|*.*DialogOptions
ofReadOnlyofPathMustExistofFileMustExist DialogTitle   Välj privat nyckelfilClickKey@AnchorsakLeftakTopakRight TabOrder TextTunnelPrivateKeyEditOnChange
DataChange    	TTabSheetSslSheetTagHelpType	htKeywordHelpKeywordui_login_tlsCaptionTLS/SSL
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxSslGroupLeft TopWidth�HeightcAnchorsakLeftakTopakRight CaptionTLS/SSL alternativTabOrder 
DesignSize�c  TLabelLabel1LeftTopWidth{HeightCaption   &Lägsta TLS/SSL-version:FocusControlMinTlsVersionCombo  TLabelLabel2LeftTop,WidthHeightCaption   &Högsta TLS/SSL-version:FocusControlMaxTlsVersionCombo  	TComboBoxMinTlsVersionComboLeft0TopWidthMHeightStylecsDropDownListAnchorsakTopakRight TabOrder OnChangeMinTlsVersionComboChangeItems.StringsSSL 2.0SSL 3.0TLS 1.0TLS 1.1TLS 1.2   	TComboBoxMaxTlsVersionComboLeft0Top'WidthMHeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChangeMaxTlsVersionComboChangeItems.StringsSSL 2.0SSL 3.0TLS 1.0TLS 1.1TLS 1.2   	TCheckBoxSslSessionReuseCheckLeftTopDWidthmHeightAnchorsakLeftakTopakRight Caption6   Å&teranvänd TLS/SSL-sessionsid för dataanslutningarTabOrderOnClick
DataChange    	TTabSheetAdvancedSheetTagHelpType	htKeywordHelpKeywordui_login_sshCaptionSSH
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxProtocolGroupLeft TopWidth�HeightWAnchorsakLeftakTopakRight Caption   Alternativ för protokollTabOrder 
DesignSize�W  TLabelLabel7LeftTop*Width� HeightCaption   Föredragen SSH-version:FocusControlSshProt1onlyButton  TRadioButtonSshProt1ButtonLeft`Top;WidthJHeightCaption&1TabOrderOnClick
DataChange  TRadioButtonSshProt2ButtonLeft� Top;WidthJHeightCaption&2TabOrderOnClick
DataChange  	TCheckBoxCompressionCheckLeftTopWidthoHeightAnchorsakLeftakTopakRight Caption   Använd &komprimeringTabOrder OnClick
DataChange  TRadioButtonSshProt1onlyButtonLeftTop;WidthJHeightCaption	End&ast 1Checked	TabOrderTabStop	OnClick
DataChange  TRadioButtonSshProt2onlyButtonLeft Top;WidthJHeightCaption	&Endast 2TabOrderOnClick
DataChange   	TGroupBoxEncryptionGroupLeft TopdWidth�Height� AnchorsakLeftakTopakRight Caption   KrypteringsinställningarTabOrder
DesignSize��   TLabelLabel8LeftTopWidth� HeightCaption$   &Riktlinjer för krypteringschiffer:FocusControlCipherListBox  TListBoxCipherListBoxLeftTop$WidthHeight[AnchorsakLeftakTopakRight DragModedmAutomatic
ItemHeightTabOrder OnClick
DataChange
OnDragDropAlgListBoxDragDrop
OnDragOverAlgListBoxDragOverOnStartDragAlgListBoxStartDrag  	TCheckBoxSsh2LegacyDESCheckLeftTop� WidthoHeightAnchorsakLeftakTopakRight Caption-   Tillåt arvsanvänding av single-&DES i SSH-2TabOrder  TButtonCipherUpButtonLeft/Top$WidthPHeightAnchorsakTopakRight Caption&UppTabOrderOnClickCipherButtonClick  TButtonCipherDownButtonLeft/TopDWidthPHeightAnchorsakTopakRight Caption&NerTabOrderOnClickCipherButtonClick    	TTabSheetKexSheetTagHelpType	htKeywordHelpKeywordui_login_kexCaption
Nyckelbyte
ImageIndex
TabVisible
DesignSize�~  	TGroupBoxKexOptionsGroupLeft TopWidth�Height� AnchorsakLeftakTopakRight Caption%   Alternativ för nyckelbytesalgoritmenTabOrder 
DesignSize��   TLabelLabel28LeftTopWidth|HeightCaption   Ri&ktlinjer för algoritmen:FocusControl
KexListBox  TListBox
KexListBoxLeftTop$WidthHeightYAnchorsakLeftakTopakRight DragModedmAutomatic
ItemHeightTabOrder OnClick
DataChange
OnDragDropAlgListBoxDragDrop
OnDragOverAlgListBoxDragOverOnStartDragAlgListBoxStartDrag  TButtonKexUpButtonLeft/Top$WidthPHeightAnchorsakTopakRight Caption&UppTabOrderOnClickKexButtonClick  TButtonKexDownButtonLeft/TopDWidthPHeightAnchorsakTopakRight Caption&NerTabOrderOnClickKexButtonClick   	TGroupBoxKexReexchangeGroupLeft Top� Width�HeightEAnchorsakLeftakTopakRight Caption(   Alternativ för kontroll av nyckelutbyteTabOrder
DesignSize�E  TLabelLabel31LeftTopWidth� HeightCaption?   Max antal minuter innan nyckeluppdatering (0 ger ingen gräns):Color	clBtnFaceFocusControlRekeyTimeEditParentColor  TLabelLabel32LeftTop,Width� HeightCaption<   Max antal data innan nyckeluppdatering (0 ger ingen gräns):Color	clBtnFaceFocusControlRekeyDataEditParentColor  TUpDownEditRekeyTimeEditLeft/TopWidthPHeight	AlignmenttaRightJustifyMaxValue       �	@AnchorsakTopakRight 	MaxLengthTabOrder OnChange
DataChange  TEditRekeyDataEditLeft/Top'WidthPHeightAnchorsakTopakRight 	MaxLength
TabOrderOnChange
DataChange    	TTabSheet	AuthSheetTagHelpType	htKeywordHelpKeywordui_login_authenticationCaptionAutentisering
ImageIndex

TabVisible
DesignSize�~  	TCheckBoxSshNoUserAuthCheckLeftTopWidth~HeightAnchorsakLeftakTopakRight Caption/   Kringgå autentisering helt och hållet (SSH-2)TabOrder OnClick
DataChange  	TGroupBoxAuthenticationGroupLeft Top Width�HeightuAnchorsakLeftakTopakRight Caption   Alternativ för autentiseringTabOrder
DesignSize�u  	TCheckBoxTryAgentCheckLeftTopWidthuHeightAnchorsakLeftakTopakRight Caption,   Försök använda autentisering med &PageantTabOrder OnClick
DataChange  	TCheckBoxAuthTISCheckLeftTop*WidthuHeightAnchorsakLeftakTopakRight Caption=   Försök använda &TIS eller Kryptokort autentisering (SSH-1)TabOrderOnClick
DataChange  	TCheckBoxAuthKICheckLeftTopAWidthuHeightAnchorsakLeftakTopakRight Caption@   Försök använda 'tagentbords&interaktiv' autentisering (SSH-2)TabOrderOnClick
DataChange  	TCheckBoxAuthKIPasswordCheckLeft TopXWidthaHeightAnchorsakLeftakTopakRight Caption)   Svara med lösenord vid första &promptenTabOrderOnClick
DataChange   	TGroupBoxAuthenticationParamsGroupLeftTop� Width�Height^AnchorsakLeftakTopakRight CaptionParametrar autentiseringTabOrder
DesignSize�^  TLabelPrivateKeyLabelLeftTop*WidthKHeightCaptionPrivat nyc&kelfilFocusControlPrivateKeyEdit  	TCheckBoxAgentFwdCheckLeftTopWidthuHeightAnchorsakLeftakTopakRight Caption   Tillåt agent-vidarebe&fordranTabOrder OnClick
DataChange  TFilenameEditPrivateKeyEditLeftTop;WidthtHeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPrivateKeyEditAfterDialogFilter8PuTTY privata nycklar (*.ppk)|*.ppk|Alla filer (*.*)|*.*DialogOptions
ofReadOnlyofPathMustExistofFileMustExist DialogTitle   Välj privat nyckelfilClickKey@AnchorsakLeftakTopakRight TabOrderTextPrivateKeyEditOnChange
DataChange   	TGroupBoxGSSAPIGroupLeft Top� Width�HeightGAnchorsakLeftakTopakRight CaptionGSSAPITabOrder
DesignSize�G  	TCheckBoxAuthGSSAPICheck3LeftTopWidthuHeightAnchorsakLeftakTopakRight Caption3   Försök använda GSSAPI/SSPI autentisering (SSH-2)TabOrder OnClickAuthGSSAPICheck3Click  	TCheckBoxGSSAPIFwdTGTCheckLeftTop*WidthuHeightAnchorsakLeftakTopakRight Caption4   Tillåt GSSAPI &vidarbefodra autentiseringsuppgifterTabOrderOnClickAuthGSSAPICheck3Click    	TTabSheet	BugsSheetTagHelpType	htKeywordHelpKeywordui_login_bugsCaptionBuggar
ImageIndex	
TabVisible
DesignSize�~  	TGroupBoxBugsGroupBoxLeft TopWidth�Height	AnchorsakLeftakTopakRight Caption   Upptäcka buggar i SSH-servrarTabOrder 
DesignSize�	  TLabelBugIgnore1LabelLeftTopWidth� HeightCaption(Stannar vid &ignore-meddelanden i SSH-1:FocusControlBugIgnore1Combo  TLabelBugPlainPW1LabelLeftTop,Width� HeightCaption*   &Vägrar all lösenordskamouflage i SSH-1:FocusControlBugPlainPW1Combo  TLabelBugRSA1LabelLeftTopDWidth� HeightCaption'Stannar vid &RSA-autentisering i SSH-1:FocusControlBugRSA1Combo  TLabelBugHMAC2LabelLeftToptWidth� HeightCaption(   Beräkningsfel av H&MAC-nycklar i SSH-2:FocusControlBugHMAC2Combo  TLabelBugDeriveKey2LabelLeftTop� Width� HeightCaption.   Beräkningsf&el av krypteringsnycklar i SSH-2:FocusControlBugDeriveKey2Combo  TLabelBugRSAPad2LabelLeftTop� Width� HeightCaption-   Kräver &utfyllnad av RSA-signaturer i SSH-2:FocusControlBugRSAPad2Combo  TLabelBugPKSessID2LabelLeftTop� Width� HeightCaption1Sessio&ns-id i SSH-2 PK autentisering missbrukas:FocusControlBugPKSessID2Combo  TLabelBugRekey2LabelLeftTop� Width� HeightCaption%   Hanterar SSH-2 nyc&kelutbyte dåligt:FocusControlBugRekey2Combo  TLabelBugMaxPkt2LabelLeftTop� Width� HeightCaption+   Ignorerar SSH-2 ma&ximum för paketstorlek:FocusControlBugMaxPkt2Combo  TLabelBugIgnore2LabelLeftTop\Width� HeightCaption(Stannar vid ignore-meddelanden i SSH-&2:FocusControlBugIgnore2Combo  	TComboBoxBugIgnore1ComboLeft@TopWidth=HeightStylecsDropDownListAnchorsakTopakRight TabOrder OnChange
DataChange  	TComboBoxBugPlainPW1ComboLeft@Top'Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugRSA1ComboLeft@Top?Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugHMAC2ComboLeft@TopoWidth=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugDeriveKey2ComboLeft@Top� Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugRSAPad2ComboLeft@Top� Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugPKSessID2ComboLeft@Top� Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugRekey2ComboLeft@Top� Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugMaxPkt2ComboLeft@Top� Width=HeightStylecsDropDownListAnchorsakTopakRight TabOrder	OnChange
DataChange  	TComboBoxBugIgnore2ComboLeft@TopWWidth=HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange     TPanel	LeftPanelLeft Top Width� Height�AlignalLeft
BevelOuterbvNoneTabOrder 
DesignSize� �  	TTreeViewNavigationTreeLeftTop	Width� Height{AnchorsakLeftakTopakRightakBottom DoubleBuffered	HideSelectionHotTrack	IndentParentDoubleBufferedReadOnly	ShowButtonsShowRootTabOrder OnChangeNavigationTreeChangeOnCollapsingNavigationTreeCollapsingItems.NodeData
�     6               ����           E n v i r o n m e n t X 6               ����            D i r e c t o r i e s X 6               ����            R e c y c l e   b i n X (               ����            S F T P X &               ����            S C P X &           ��������            F T P X 4               ����           C o n n e c t i o n X *               ����            P r o x y X ,               ����            T u n n e l X &               ����           S S H X 8               ����            K e x   e x c h a n g e X <               ����            A u t h e n t i c a t i o n X (               ����            B u g s X     TButtonOKBtnLeft3Top�WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft�Top�WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeft�Top�WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TButtonColorButtonLeftTop�WidthRHeightAnchorsakLeftakBottom Caption   &FärgTabOrderOnClickColorButtonClick  
TImageListColorImageListAllocByLefttTop�Bitmap
&  IL  P   �������������BM6       6   (   @                                                                                                                                                                                                                                                                                                                K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5                                                                                                                                                                                                                                         K?5 K?5 K?5 K?5                                                                                                                                                                                                                             dYQ K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 bXO                                                                                                                                                                                                         K?5 s`R s`R s`R s`R s`R s`R s`R s`R s`R s`R s`R s`R K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         bXO K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 bXO                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     BM>       >   (   @            �                       ��� ��      �      �?      �      �      �      �      �      �      �      �      �      �      �      ��      ��                                  TPF0TSymlinkDialogSymlinkDialogLeft�Top� HelpType	htKeywordHelpKeyword
ui_symlinkBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSymlinkDialogClientHeight� ClientWidth�Color	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenterOnShowFormShow
DesignSize��  PixelsPerInch`
TextHeight 	TGroupBoxSymlinkGroupLeftTopWidth|Height� AnchorsakLeftakTopakRightakBottom TabOrder 
DesignSize|�   TLabelFileNameLabelLeftTopWidthSHeightCaption   &Länk/genväg fil:FocusControlFileNameEdit  TLabelLabel1LeftTop@WidthgHeightCaption   &Pekar länk/genväg till:FocusControlPointToEdit  TEditFileNameEditLeftTop WidthfHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeControlChange  TEditPointToEditLeftTopPWidthfHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChange  	TCheckBoxSymbolicCheckLeftTopmWidth� HeightCaption   Sy&mbolisk länkTabOrderOnClickControlChange   TButtonOkButtonLeft� Top� WidthKHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top� WidthKHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeft8Top� WidthKHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick     TPF0TSynchronizeChecklistDialogSynchronizeChecklistDialogLeft4Top� HelpType	htKeywordHelpKeywordui_synchronize_checklistBorderIconsbiSystemMenu
biMaximizebiHelp Caption   Checklist för synkroniseringClientHeight�ClientWidth�Color	clBtnFaceConstraints.MinHeight^Constraints.MinWidth|
ParentFont		Icon.Data
~           h     (                 @                           [��![��![��![��![��![��![��![��![��![��![�� [��                ![��+f��+f��+f��+f��+f��+f��+f��+f��+f��+f��![��                ![��l�����������������������������������,h��![��                ![��m�����������������������������������-i��![��                ![��n�����������{w����pm��������������.k��![��                ![��o�����������54��������������������/l��![��                ![��p�������������������qn��qn����������0n��![��                ![��q���������������������������������1p��![��                ![��r�����������������������qo��qo������2q��![��                ![��s���������������������������������3r��![��                ![��t�����������������������������������4t��![��                ![��t�����������������������������������4t��![��                ![������t���SPP�SPP�SPP�SPP�SPP�SPP�t���4t��![��                !\��![��![��������������������������![��![��!\��                            SPP�SPP�SQQ�SQQ�SPP�SPP�                                            TOOjSPP�SPP�TOOj                        �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �?  
KeyPreview	OldCreateOrder	PositionpoOwnerFormCenterOnShowFormShowPixelsPerInch`
TextHeight TPanelPanelLeft;Top Width|Height�AlignalRight
BevelOuterbvNoneTabOrder
DesignSize|�  TButtonOkButtonLeftTopWidthlHeightAnchorsakLeftakTopakRight CaptionOKDefault	ModalResultTabOrder   TButtonCancelButtonLeftTop(WidthlHeightAnchorsakLeftakTopakRight Cancel	CaptionAvbrytModalResultTabOrder  TButtonCheckAllButtonLeftTop� WidthlHeightAnchorsakLeftakTopakRight CaptionMarkera &allaTabOrderOnClickCheckAllButtonClick  TButtonUncheckAllButtonLeftTop� WidthlHeightAnchorsakLeftakTopakRight CaptionAvmarkera a&llaTabOrderOnClickCheckAllButtonClick  TButtonCheckButtonTagLeftTopvWidthlHeightAnchorsakLeftakTopakRight CaptionMarkeraTabOrderOnClickCheckButtonClick  TButtonUncheckButtonLeftTop� WidthlHeightAnchorsakLeftakTopakRight Caption	AvmarkeraTabOrderOnClickCheckButtonClick  TButton
HelpButtonLeftTopHWidthlHeightAnchorsakLeftakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick  TButtonCustomCommandsButtonTagLeftTopWidthlHeightAnchorsakLeftakTopakRight CaptionEgna ko&mmandonTabOrderOnClickCustomCommandsButtonClick   TIEListViewListViewLeft Top Width;Height�AlignalClient
Checkboxes	FullDrag	HideSelectionReadOnly		RowSelect		PopupMenuListViewPopupMenuTabOrder 	ViewStylevsReportOnChangeListViewChange
OnChangingListViewChanging
NortonLikenlOffColumnsCaptionNamn CaptionLokal katalogWidthd 	AlignmenttaRightJustifyCaptionStorlekWidthF Caption   ÄndradWidthP MaxWidthMinWidthWidth Caption   FjärrkatalogWidthd 	AlignmenttaRightJustifyCaptionStorlekWidthF Caption   ÄndradWidthP  OnAdvancedCustomDrawSubItem!ListViewAdvancedCustomDrawSubItem	OnCompareListViewCompareOnContextPopupListViewContextPopupOnSelectItemListViewSelectItemOnSecondaryColumnHeaderListViewSecondaryColumnHeader  
TStatusBar	StatusBarLeft Top�Width�HeightHint9   Klicka för att markera alla åtgärder av den här typenPanelsStylepsOwnerDrawText'   Fullständiga synkroniseringsåtgärderWidth_ StylepsOwnerDrawTextNya lokala filerWidth_ StylepsOwnerDrawText   Nya fjärrfilerWidth_ StylepsOwnerDrawTextUppdaterade lokala filerWidth_ StylepsOwnerDrawText   Uppdaterade fjärrfilerWidth_ StylepsOwnerDrawText   Gamla fjärrfilerWidth_ StylepsOwnerDrawTextGamla lokala filerWidth_ Width2  ParentShowHintShowHint	OnMouseDownStatusBarMouseDownOnMouseMoveStatusBarMouseMoveOnDrawPanelStatusBarDrawPanel  TPngImageListActionImages	PngImages
BackgroundclWindowName2Total actions counter on synchronization checklistPngImage.Data
x  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATx�c���?0222 ��,F�� ����7���,ׇ̀����@*(�Q�P��oذ6�3c�3�g����71`�:� F�#��٢���79��Ǘ���c5�7I��¡���eH_r�� ��`�.|`K�~$=:�j|�g7�����f�8�1H�c���+�-�f~'�2���bx��v�B��1�p��L�w3�6cx��=v�D���}��9���bb{��{����"����d���a`f�P]�7h���ڔ��ۏ����c��f�9���ɦ����0�fp>x��CT�n�)Ç���`��� �N|���͝� àی���j�O>c7��Ǉ�ߣ��������p��U&�?}�n���7�{/ބt�ژ�������b |��Ӏ1�G��1�?��cK�[�� �w��yhM    IEND�B`� 
BackgroundclWindowNameNew local files indicatorPngImage.Data
S  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   �IDATx�c���?%�q@�B�v���������N�B���4n\����Y��. �.th���̑���l���p�tb����ٳ�>����O�,F����8ؖG�^2<�|�Sd 33��˗�=��*���z�P�%1�^�8)�ƁO�n  䳚w�]��    IEND�B`� 
BackgroundclWindowNameNew remote files indicatorPngImage.Data
X  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   �IDATx�c���?%�q�̑��������*�;�d�B�p<3�4%��W�2<�|�H�RR\l�?�������2�g��pt�I���B���؀=z�a�;[t1F�v�c�
ʖ��:��~c���� ��93q�M�N��*F��� T|��
��@1Kt1���h��8�  �e�dI���    IEND�B`� 
BackgroundclWindowNameModified local files indicatorPngImage.Data
R  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   �IDATx�c���?%�q@��Y����32
0������u������@^����g���������B�@��@���H��϶8����0|��̭���~_��Û2�X�_���q��`��`����p��C��O����G��@���;���%1�^�8)�ƁO�n  Ͳ��<�s�    IEND�B`� 
BackgroundclWindowNameModified remote files indicatorPngImage.Data
R  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�   �IDATx�c���?%�q�̙�ã���i��i�?;�d�L^�xff�i:b"\_�bH����(fJIq1|�<���3�XQ������7����{����P�]�蘜�����<�o�?}A6�X�_���Q� �^8
TgR���>[��Q�G����7  �P>�֠    IEND�B`� 
BackgroundclWindowNameObsolete local files indicatorPngImage.Data
v  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڥ�KLSQ��>z���ii�
mx*A�+$l\FcܰacK01х_�.\ibԴcdc4���Mc"�GRT�h�1��}Ж>���� .<�33����?���P*��(��[��~��G��l�|���g2��&J�GNJ҄�3����/܍��ӡ��J�v{Dq`mq?B�<�!�k�A��
����G�\�oF��8+ �$ax$�K�f��HҐZ|���h�
�V;��Z�0��gA�� >tحG[v6 I��(�Hp<���S:]�ٗ;ꪜ��
�����\0�7��..��1Eq1�߳!Ե��X��eA�W�2�������R�/��td0�{%)��W�2 �@�TTt����X��q��ߢ1x?=�����Gԧ�(?�/��W�U���鴻2M0<%�y$i���	 uq}����Z��n&��O?��Ц��)�t�ճ���2�'݅��6��9�"��4�N--�� >��|�\k%;6Wr9x�S�3{l%�|L����$u� ���-躉a��E8�ƴ�������Mڄ�y3"f�8�d���<!����R0�r��h��������(��Wo�����wRp�v�N�R)�f�>�֞_ s'xp�r_�y�0\%�k��3�k �����H��\�8��G�:�,In�W��n�����
%�>%����u�&��������������'�zn�K��    IEND�B`� 
BackgroundclWindowNameObsolete remote files indicatorPngImage.Data
v  �PNG

   IHDR         ��a   	pHYs  �  ��+  
OiCCPPhotoshop ICC profile  xڝSgTS�=���BK���KoR RB���&*!	J�!��Q�EEȠ�����Q,�
��!���������{�kּ������>�����H3Q5��B�������.@�
$p �d!s�# �~<<+"�� x� �M��0���B�\���t�8K� @z�B� @F���&S � `�cb� P- `'�� ����{ [�!��  e�D h; ��V�E X0 fK�9 �- 0IWfH �� ���  0Q��) { `�##x �� F�W<�+��*  x��<�$9E�[-qWW.(�I+6aa�@.�y�2�4���  ������x����6��_-��"bb���ϫp@  �t~��,/��;�m��%�h^�u��f�@� ���W�p�~<<E���������J�B[a�W}�g�_�W�l�~<�����$�2]�G�����L�ϒ	�b��G�����"�Ib�X*�Qq�D���2�"�B�)�%��d��,�>�5 �j>{�-�]c�K'Xt���  �o��(�h���w��?�G�% �fI�q  ^D$.Tʳ?�  D��*�A��,�����`6�B$��BB
d�r`)��B(�Ͱ*`/�@4�Qh��p.�U�=p�a��(��	A�a!ڈb�X#����!�H�$ ɈQ"K�5H1R�T UH�=r9�\F��;� 2����G1���Q=��C��7�F��dt1�����r�=�6��Ыhڏ>C�0��3�l0.��B�8,	�c˱"����V����cϱw�E�	6wB aAHXLXN�H� $4�	7	�Q�'"��K�&���b21�XH,#��/{�C�7$�C2'��I��T��F�nR#�,��4H#���dk�9�, +ȅ����3��!�[
�b@q��S�(R�jJ��4�e�2AU��Rݨ�T5�ZB���R�Q��4u�9̓IK�����hh�i��t�ݕN��W���G���w��ǈg(�gw��L�Ӌ�T071���oUX*�*|��
�J�&�*/T����ުU�U�T��^S}�FU3S�	Ԗ�U��P�SSg�;���g�oT?�~Y��Y�L�OC�Q��_�� c�x,!k��u�5�&���|v*�����=���9C3J3W�R�f?�q��tN	�(���~���)�)�4L�1e\k����X�H�Q�G�6����E�Y��A�J'\'Gg����S�Sݧ
�M=:��.�k���Dw�n��^��Lo��y���}/�T�m���GX�$��<�5qo</���QC]�@C�a�a�ᄑ��<��F�F�i�\�$�m�mƣ&&!&KM�M�RM��)�;L;L���͢�֙5�=1�2��כ߷`ZxZ,����eI��Z�Yn�Z9Y�XUZ]�F���%ֻ�����N�N���gð�ɶ�����ۮ�m�}agbg�Ů��}�}��=���Z~s�r:V:ޚΜ�?}����/gX���3��)�i�S��Ggg�s�󈋉K��.�>.���Ƚ�Jt�q]�z��������ۯ�6�i�ܟ�4�)�Y3s���C�Q��?��0k߬~OCO�g��#/c/�W�װ��w��a�>�>r��>�<7�2�Y_�7��ȷ�O�o�_��C#�d�z�� ��%g��A�[��z|!��?:�e����A���AA�������!h�쐭!��Α�i�P~���a�a��~'���W�?�p�X�1�5w��Cs�D�D�Dޛg1O9�-J5*>�.j<�7�4�?�.fY��X�XIlK9.*�6nl��������{�/�]py�����.,:�@L�N8��A*��%�w%�
y��g"/�6ш�C\*N�H*Mz�쑼5y$�3�,幄'���LLݛ:��v m2=:�1����qB�!M��g�g�fvˬe����n��/��k���Y-
�B��TZ(�*�geWf�͉�9���+��̳�ې7�����ᒶ��KW-X潬j9�<qy�
�+�V�<���*m�O��W��~�&zMk�^�ʂ��k�U
�}����]OX/Yߵa���>������(�x��oʿ�ܔ���Ĺd�f�f���-�[����n�ڴ�V����E�/��(ۻ��C���<��e����;?T�T�T�T6��ݵa��n��{��4���[���>ɾ�UUM�f�e�I���?�������m]�Nmq����#�׹���=TR��+�G�����w-6U����#pDy���	��:�v�{���vg/jB��F�S��[b[�O�>����z�G��4<YyJ�T�i��ӓg�ό���}~.��`ۢ�{�c��jo�t��E���;�;�\�t���W�W��:_m�t�<���Oǻ�����\k��z��{f���7����y���՞9=ݽ�zo������~r'��˻�w'O�_�@�A�C݇�?[�����j�w����G��������C���ˆ��8>99�?r����C�d�&����ˮ/~�����јѡ�򗓿m|������������x31^�V���w�w��O�| (�h���SЧ��������c3-�  �IDATxڥ�KLSQ��>z���ii�
mx*A�+$l\FcܰacK01х_�.\ibԴcdc4���Mc"�GRT�h�1��}Ж>���� .<�33����?���P*��(��[��~��G��l�|���g2��&J�GNJ҄�3����/܍��ӡ��J�v{Dq`mq?B�<�!�k�A��
����G�\�oF��8+ �$ax$�K�f��HҐZ|���h�
�V;��Z�0��gA�� >tحG[v6 I��(�Hp<���S:]�ٗ;ꪜ��
�����\0�7��..��1Eq1�߳!Ե��X��eA�W�2�������R�/��td0�{%)��W�2 �@�TTt����X��q��ߢ1x?=�����Gԧ�(?�/��W�U���鴻2M0<%�y$i���	 uq}����Z��n&��O?��Ц��)�t�ճ���2�'݅��6��9�"��4�N--�� >��|�\k%;6Wr9x�S�3{l%�|L����$u� ���-躉a��E8�ƴ�������Mڄ�y3"f�8�d���<!����R0�r��h��������(��Wo�����wRp�v�N�R)�f�>�֞_ s'xp�r_�y�0\%�k��3�k �����H��\�8��G�:�,In�W��n�����
%�>%����u�&��������������'�zn�K��    IEND�B`�  LefthTophBitmap
      
TPopupMenuListViewPopupMenuLefthTopH 	TMenuItem	CheckItemTagCaption&MarkeraOnClickCheckButtonClick  	TMenuItemUncheckItemCaption
&AvmarkeraOnClickCheckButtonClick  	TMenuItemN1Caption-  	TMenuItemSelectAllItemCaption&Markera allaShortCutA@OnClickSelectAllItemClick   TTimerUpdateTimerEnabledIntervaldOnTimerUpdateTimerTimerLefthTop(  
TImageListArrowImagesLeft�TophBitmap
&  IL     �������������BM6       6   (   @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ��� ��� ��� ��� ��� ��� ��� ���                                             ��� ���                                                                                                                                                                             ���                         ���                                         ���         ���                                                                                                                                                                             ���                 ���                                             ���         ���                                                                                                                                                                             ���                 ���                                         ���                 ���                                                                                                                                                                             ���         ���                                             ���                 ���                                                                                                                                                                             ���         ���                                         ���                         ���                                                                                                                                                                             ��� ���                                             ��� ��� ��� ��� ��� ��� ��� ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 BM>       >   (   @            �                       ��� ����    ����    ����    ����    ����    ��    ����    ����    ����    ����    ����    ��    ����    ����    ����    ����                              TPF0TSynchronizeDialogSynchronizeDialogLeftoTop� HelpType	htKeywordHelpKeywordui_keepuptodateBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption"Keep remote directory up to date XClientHeight�ClientWidth�Color	clBtnFace
ParentFont	
KeyPreview	OldCreateOrderPositionpoOwnerFormCenterOnCloseQueryFormCloseQuery	OnKeyDownFormKeyDownOnShowFormShow
DesignSize�� PixelsPerInch`
TextHeight 	TGroupBoxDirectoriesGroupLeftTopWidth�HeightwAnchorsakLeftakTopakRight Caption	KatalogerTabOrder 
DesignSize�w  TLabelLocalDirectoryLabelLeft1TopWidth� HeightAnchorsakLeftakTopakRight Caption.   Be&vaka förändringar i den lokala katalogen:FocusControlLocalDirectoryEdit  TLabelRemoteDirectoryLabelLeft1TopDWidthHeightAnchorsakLeftakTopakRight Caption6   ... och inför dessa &automatiskt på fjärrkatalogen:FocusControlRemoteDirectoryEdit  TImageImageLeftTopWidth Height AutoSize	Picture.Data
Z  	TPngImage�PNG

   IHDR           szz�   	pHYs  �  ��o�d  IDATx�ŗkLU��wf��Ky����Zb�����Fi+���
M��hk|4i��4��"јچ���Š_L�"���H
m
��,�²��Lمe����x6�{f��=�{���%���x����|Fx���<�?/*x�?��"y�nq�ż='���.\��#�77�w��A\V����*���84ph镜�'[�bx�xk�6�6�c��;q����}�c����1J�^��?1<�z�G:��)���X����8˭2� ��V�5�	�՝wP{��^�(�J�
J��#p�ݰZ�1t��9γ��)�2��f�h�[~A_�����Bg}���l�����\����BJ	#}�9Cw����Mdef"9!�ϟ	�V�Rp�ӆ�ڝU�!UH1iq��%�B��!>��H�iJȊB��O�;��F`��y^i��f��G2�,��J�
�E5;�:8�G��d��^�Z+��R?��g�8����[�6�n�LB��Ix>-�w�B���/��Zs@��U�[��Ѩ�~K#���k� �U~�� =V^m��1(I���k8����a�����%�%̪	jN�x���&�7����P�>�m��\�I�O�K�0{��GO	(ػ0����`����3+3C�8. ��`����9@ø ��t��� @�j��tE����@8�ؐ�a��R�0��Ң��l�}�{����^�����'�"�ź�g�)����磑���������������WĚ��҆��&�a��މ��� �cW���.7�r����0����3�I BU�93�qfp �~h��iP�y/��q��=6���Z/���s/AW��t�.߬��h��]�-<�?��jm�S��s&�Q;��O�C���`J=� �o�0�z����R�Un��>�l��0C=�֛�Ryn���FB�f^ �z�l�[wo6���o ���V���.�~���Kn;C�[0�퀂�\�B�'�!-�W=� �6o��7U���8
34:���qL`<5aK��{<J`��Xdj&4 ��� O�apЄ��kX���h=��������8�.\���<S���� �y|%���y��Lxf�\�/Y��2�hW��ä�	��	#l$�ܩĚ=jH���i^���j��h��{���&�!��'x�v�Z�;�<E���9IN(���|�y��pD��c	���l�jr$����z�p���R}pт��
���Aڿ�D�?��    IEND�B`�  THistoryComboBoxRemoteDirectoryEditLeft1TopTWidthiHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeControlChange  THistoryComboBoxLocalDirectoryEditLeft1Top#WidthHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder TextLocalDirectoryEditOnChangeControlChange  TButtonLocalDirectoryBrowseButtonLeftOTop!WidthKHeightAnchorsakTopakRight Caption   &Bläddra...TabOrderOnClickLocalDirectoryBrowseButtonClick   TButton
StopButtonLeft� Top WidthJHeightAnchorsakTopakRight Caption&StoppTabOrderOnClickStopButtonClick  TButtonCancelButtonLeftTop WidthJHeightAnchorsakTopakRight Cancel	Caption   StängModalResultTabOrder  	TGroupBoxOptionsGroupLeftTop� Width�Height_AnchorsakLeftakTopakRight Caption   Alternativ för synkroniseringTabOrder
DesignSize�_  	TCheckBoxSynchronizeDeleteCheckLeftTopWidth� HeightCaption&Ta bort filerTabOrder OnClickControlChange  	TCheckBoxSaveSettingsCheckLeftTopDWidth� HeightCaption*   Använd &samma inställningar nästa gångTabOrderOnClickControlChange  	TCheckBoxSynchronizeExistingOnlyCheckLeft� TopWidth� HeightAnchorsakLeftakTopakRight CaptionBara &existerande filerTabOrderOnClickControlChange  	TCheckBoxSynchronizeRecursiveCheckLeftTop,Width� HeightCaption&Uppdatera underkatalogerTabOrderOnClickControlChange  TGrayedCheckBoxSynchronizeSynchronizeCheckLeft� TopDWidth� HeightAllowGrayed	AnchorsakLeftakTopakRight CaptionSynkronisera vid s&tartTabOrderOnClickControlChange  	TCheckBoxSynchronizeSelectedOnlyCheckLeft� Top,Width� HeightCaption&Bara markerade filerTabOrderOnClickControlChange   TButtonStartButtonLeft� Top WidthJHeightAnchorsakTopakRight Caption&StartDefault	TabOrderOnClickStartButtonClick  TButtonMinimizeButtonLeftTop WidthJHeightAnchorsakTopakRight Caption	&MinimeraTabOrderOnClickMinimizeButtonClick  TButtonTransferSettingsButtonLeftTop Width� HeightCaption   Över&föringsinställningarTabOrderOnClickTransferSettingsButtonClickOnDropDownClick#TransferSettingsButtonDropDownClick  	TGroupBoxCopyParamGroupLeftTop� Width�Height2AnchorsakLeftakTopakRight Caption   ÖverföringsinställningarTabOrderOnClickCopyParamGroupClickOnContextPopupCopyParamGroupContextPopup
DesignSize�2  TLabelCopyParamLabelLeftTopWidth�HeightAnchorsakLeftakTopakRightakBottom AutoSizeCaptionCopyParamLabelWordWrap	OnClickCopyParamGroupClick   TButton
HelpButtonLeftaTop WidthKHeightAnchorsakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick  TPanelLogPanelLeft TopAWidth�HeightdAlignalBottom
BevelOuterbvNoneTabOrder	
DesignSize�d  	TListViewLogViewLeftTopWidth�HeightZAnchorsakLeftakTopakRightakBottom ColumnsWidth�	WidthType�  Width�	WidthType�   DoubleBuffered	ReadOnly		RowSelect	ParentDoubleBufferedShowColumnHeadersTabOrder 	ViewStylevsReport	OnKeyDownLogViewKeyDown    TPF0TSynchronizeProgressFormSynchronizeProgressFormLeftOTopBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSynchronization XClientHeightClientWidth~Color	clBtnFace
ParentFont	OldCreateOrderPositionpoOwnerFormCenter
DesignSize~ PixelsPerInch`
TextHeight TLabelLabel1LeftTop	WidthHeightCaptionLokal:  TLabelLabel2LeftTopWidth)HeightCaption   Fjärr:  
TPathLabelRemoteDirectoryLabelLefteTopWidthHeightUnixPath	IndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  
TPathLabelLocalDirectoryLabelLeftdTop	WidthHeightIndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TLabelStartTimeLabelLeftdTop1WidthQHeightAutoSizeCaption00:00:00  TLabelLabel4LeftTop1Width3HeightCaptionStartad:  TLabelLabel3LeftTopEWidthBHeightCaption   Förfluten tid:  TLabelTimeElapsedLabelLeftdTopEWidthOHeightAutoSizeCaption00:00:00  TButtonCancelButtonLeft� Top^WidthIHeightAnchorsakRightakBottom CaptionAvbrytTabOrder OnClickCancelButtonClick  TButtonMinimizeButtonLeft-Top^WidthIHeightAnchorsakRightakBottom Caption	&MinimeraTabOrderOnClickMinimizeButtonClick  TTimerUpdateTimerEnabledOnTimerUpdateTimerTimerLeft)TopY         @   4        �      D4   V S _ V E R S I O N _ I N F O     ���   =                                     �    S t r i n g F i l e I n f o   ~    0 4 1 D f d e 9   >   C o m p a n y N a m e     M a r t i n   P r i k r y l     n #  F i l e D e s c r i p t i o n     S w e d i s h   t r a n s l a t i o n   o f   W i n S C P   ( S V )     *   F i l e V e r s i o n     1 . 6 1     � 3  L e g a l C o p y r i g h t   ( c )   2 0 0 3 - 2 0 1 4   A n d r e a s   P e t t e r s s o n   a n d   R e n � �   F i c h t e r     < 
  O r i g i n a l F i l e n a m e   W i n S C P . s v   4   P r o d u c t V e r s i o n   5 . 5 . 4 . 0   6   W W W     h t t p : / / w i n s c p . n e t /     (   L a n g N a m e   S w e d i s h   .   P r o d u c t N a m e     W i n S C P     D     V a r F i l e I n f o     $    T r a n s l a t i o n     ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        